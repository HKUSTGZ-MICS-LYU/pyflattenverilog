// Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:1
module b19(clock, reset, bs, na, hold, in1, in2, in3, ris);
    input clock;
    input reset;
    input bs;
    input na;
    input hold;
    input [10:0] in1;
    input [10:0] in2;
    input [19:0] in3;
    output [29:0] ris;

    reg P1_P1_P1_ADS_n = 1'b0;
    reg [29:0] P1_P1_P1_Address = 30'b0;
    reg [3:0] P1_P1_P1_BE_n = 4'b0;
    reg P1_P1_P1_BS16_n = 1'b0;
    reg [3:0] P1_P1_P1_ByteEnable = 4'b0;
    reg P1_P1_P1_CLOCK = 1'b0;
    reg P1_P1_P1_CodeFetch = 1'b0;
    reg P1_P1_P1_D_C_n = 1'b0;
    reg signed [31:0] P1_P1_P1_DataWidth = 32'b0;
    reg [31:0] P1_P1_P1_Datai = 32'b0;
    reg signed [31:0] P1_P1_P1_Datao = 32'b0;
    reg signed [31:0] P1_P1_P1_EAX = 32'b0;
    reg signed [31:0] P1_P1_P1_EBX = 32'b0;
    reg P1_P1_P1_Extended = 1'b0;
    reg P1_P1_P1_Flush = 1'b0;
    reg P1_P1_P1_HOLD = 1'b0;
    reg signed [31:0] P1_P1_P1_InstAddrPointer = 32'b0;
    reg [7:0] P1_P1_P1_InstQueue [15:0];
    reg [4:0] P1_P1_P1_InstQueueRd_Addr = 5'b0;
    reg [4:0] P1_P1_P1_InstQueueWr_Addr = 5'b0;
    reg P1_P1_P1_M_IO_n = 1'b0;
    reg P1_P1_P1_MemoryFetch = 1'b0;
    reg P1_P1_P1_More = 1'b0;
    reg P1_P1_P1_NA_n = 1'b0;
    reg P1_P1_P1_NonAligned = 1'b0;
    reg signed [31:0] P1_P1_P1_PhyAddrPointer = 32'b0;
    reg P1_P1_P1_READY_n = 1'b0;
    reg P1_P1_P1_RESET = 1'b0;
    reg P1_P1_P1_ReadRequest = 1'b0;
    reg P1_P1_P1_RequestPending = 1'b0;
    reg [2:0] P1_P1_P1_State = 3'b0;
    reg [3:0] P1_P1_P1_State2 = 4'b0;
    reg P1_P1_P1_StateBS16 = 1'b0;
    reg P1_P1_P1_StateNA = 1'b0;
    reg P1_P1_P1_W_R_n = 1'b0;
    reg signed [31:0] P1_P1_P1_fWord = 32'b0;
    reg [15:0] P1_P1_P1_lWord = 16'b0;
    reg signed [31:0] P1_P1_P1_rEIP = 32'b0;
    reg [14:0] P1_P1_P1_uWord = 15'b0;
    reg P1_P1_P2_ADS_n = 1'b0;
    reg [29:0] P1_P1_P2_Address = 30'b0;
    reg [3:0] P1_P1_P2_BE_n = 4'b0;
    reg P1_P1_P2_BS16_n = 1'b0;
    reg [3:0] P1_P1_P2_ByteEnable = 4'b0;
    reg P1_P1_P2_CLOCK = 1'b0;
    reg P1_P1_P2_CodeFetch = 1'b0;
    reg P1_P1_P2_D_C_n = 1'b0;
    reg signed [31:0] P1_P1_P2_DataWidth = 32'b0;
    reg [31:0] P1_P1_P2_Datai = 32'b0;
    reg signed [31:0] P1_P1_P2_Datao = 32'b0;
    reg signed [31:0] P1_P1_P2_EAX = 32'b0;
    reg signed [31:0] P1_P1_P2_EBX = 32'b0;
    reg P1_P1_P2_Extended = 1'b0;
    reg P1_P1_P2_Flush = 1'b0;
    reg P1_P1_P2_HOLD = 1'b0;
    reg signed [31:0] P1_P1_P2_InstAddrPointer = 32'b0;
    reg [7:0] P1_P1_P2_InstQueue [15:0];
    reg [4:0] P1_P1_P2_InstQueueRd_Addr = 5'b0;
    reg [4:0] P1_P1_P2_InstQueueWr_Addr = 5'b0;
    reg P1_P1_P2_M_IO_n = 1'b0;
    reg P1_P1_P2_MemoryFetch = 1'b0;
    reg P1_P1_P2_More = 1'b0;
    reg P1_P1_P2_NA_n = 1'b0;
    reg P1_P1_P2_NonAligned = 1'b0;
    reg signed [31:0] P1_P1_P2_PhyAddrPointer = 32'b0;
    reg P1_P1_P2_READY_n = 1'b0;
    reg P1_P1_P2_RESET = 1'b0;
    reg P1_P1_P2_ReadRequest = 1'b0;
    reg P1_P1_P2_RequestPending = 1'b0;
    reg [2:0] P1_P1_P2_State = 3'b0;
    reg [3:0] P1_P1_P2_State2 = 4'b0;
    reg P1_P1_P2_StateBS16 = 1'b0;
    reg P1_P1_P2_StateNA = 1'b0;
    reg P1_P1_P2_W_R_n = 1'b0;
    reg signed [31:0] P1_P1_P2_fWord = 32'b0;
    reg [15:0] P1_P1_P2_lWord = 16'b0;
    reg signed [31:0] P1_P1_P2_rEIP = 32'b0;
    reg [14:0] P1_P1_P2_uWord = 15'b0;
    reg P1_P1_P3_ADS_n = 1'b0;
    reg [29:0] P1_P1_P3_Address = 30'b0;
    reg [3:0] P1_P1_P3_BE_n = 4'b0;
    reg P1_P1_P3_BS16_n = 1'b0;
    reg [3:0] P1_P1_P3_ByteEnable = 4'b0;
    reg P1_P1_P3_CLOCK = 1'b0;
    reg P1_P1_P3_CodeFetch = 1'b0;
    reg P1_P1_P3_D_C_n = 1'b0;
    reg signed [31:0] P1_P1_P3_DataWidth = 32'b0;
    reg [31:0] P1_P1_P3_Datai = 32'b0;
    reg signed [31:0] P1_P1_P3_Datao = 32'b0;
    reg signed [31:0] P1_P1_P3_EAX = 32'b0;
    reg signed [31:0] P1_P1_P3_EBX = 32'b0;
    reg P1_P1_P3_Extended = 1'b0;
    reg P1_P1_P3_Flush = 1'b0;
    reg P1_P1_P3_HOLD = 1'b0;
    reg signed [31:0] P1_P1_P3_InstAddrPointer = 32'b0;
    reg [7:0] P1_P1_P3_InstQueue [15:0];
    reg [4:0] P1_P1_P3_InstQueueRd_Addr = 5'b0;
    reg [4:0] P1_P1_P3_InstQueueWr_Addr = 5'b0;
    reg P1_P1_P3_M_IO_n = 1'b0;
    reg P1_P1_P3_MemoryFetch = 1'b0;
    reg P1_P1_P3_More = 1'b0;
    reg P1_P1_P3_NA_n = 1'b0;
    reg P1_P1_P3_NonAligned = 1'b0;
    reg signed [31:0] P1_P1_P3_PhyAddrPointer = 32'b0;
    reg P1_P1_P3_READY_n = 1'b0;
    reg P1_P1_P3_RESET = 1'b0;
    reg P1_P1_P3_ReadRequest = 1'b0;
    reg P1_P1_P3_RequestPending = 1'b0;
    reg [2:0] P1_P1_P3_State = 3'b0;
    reg [3:0] P1_P1_P3_State2 = 4'b0;
    reg P1_P1_P3_StateBS16 = 1'b0;
    reg P1_P1_P3_StateNA = 1'b0;
    reg P1_P1_P3_W_R_n = 1'b0;
    reg signed [31:0] P1_P1_P3_fWord = 32'b0;
    reg [15:0] P1_P1_P3_lWord = 16'b0;
    reg signed [31:0] P1_P1_P3_rEIP = 32'b0;
    reg [14:0] P1_P1_P3_uWord = 15'b0;
    reg [29:0] P1_P1_addr1 = 30'b0;
    reg [29:0] P1_P1_addr2 = 30'b0;
    reg [29:0] P1_P1_addr3 = 30'b0;
    reg [29:0] P1_P1_address1 = 30'b0;
    reg [29:0] P1_P1_address2 = 30'b0;
    reg P1_P1_ads1 = 1'b0;
    reg P1_P1_ads2 = 1'b0;
    reg P1_P1_ads3 = 1'b0;
    reg P1_P1_ast1 = 1'b0;
    reg P1_P1_ast2 = 1'b0;
    reg [3:0] P1_P1_be1 = 4'b0;
    reg [3:0] P1_P1_be2 = 4'b0;
    reg [3:0] P1_P1_be3 = 4'b0;
    reg P1_P1_bs16 = 1'b0;
    reg signed [31:0] P1_P1_buf1 = 32'b0;
    reg signed [31:0] P1_P1_buf2 = 32'b0;
    reg P1_P1_clock = 1'b0;
    reg [31:0] P1_P1_datai = 32'b0;
    reg signed [31:0] P1_P1_datao = 32'b0;
    reg P1_P1_dc = 1'b0;
    reg P1_P1_dc1 = 1'b0;
    reg P1_P1_dc2 = 1'b0;
    reg P1_P1_dc3 = 1'b0;
    reg signed [31:0] P1_P1_di1 = 32'b0;
    reg signed [31:0] P1_P1_di2 = 32'b0;
    reg signed [31:0] P1_P1_di3 = 32'b0;
    reg [31:0] P1_P1_do1 = 32'b0;
    reg [31:0] P1_P1_do2 = 32'b0;
    reg [31:0] P1_P1_do3 = 32'b0;
    reg P1_P1_hold = 1'b0;
    reg P1_P1_mio = 1'b0;
    reg P1_P1_mio1 = 1'b0;
    reg P1_P1_mio2 = 1'b0;
    reg P1_P1_mio3 = 1'b0;
    reg P1_P1_na = 1'b0;
    reg P1_P1_rdy1 = 1'b0;
    reg P1_P1_rdy2 = 1'b0;
    reg P1_P1_rdy3 = 1'b0;
    reg P1_P1_ready1 = 1'b0;
    reg P1_P1_ready11 = 1'b0;
    reg P1_P1_ready12 = 1'b0;
    reg P1_P1_ready2 = 1'b0;
    reg P1_P1_ready21 = 1'b0;
    reg P1_P1_ready22 = 1'b0;
    reg P1_P1_reset = 1'b0;
    reg P1_P1_wr = 1'b0;
    reg P1_P1_wr1 = 1'b0;
    reg P1_P1_wr2 = 1'b0;
    reg P1_P1_wr3 = 1'b0;
    reg P1_P2_P1_ADS_n = 1'b0;
    reg [29:0] P1_P2_P1_Address = 30'b0;
    reg [3:0] P1_P2_P1_BE_n = 4'b0;
    reg P1_P2_P1_BS16_n = 1'b0;
    reg [3:0] P1_P2_P1_ByteEnable = 4'b0;
    reg P1_P2_P1_CLOCK = 1'b0;
    reg P1_P2_P1_CodeFetch = 1'b0;
    reg P1_P2_P1_D_C_n = 1'b0;
    reg signed [31:0] P1_P2_P1_DataWidth = 32'b0;
    reg [31:0] P1_P2_P1_Datai = 32'b0;
    reg signed [31:0] P1_P2_P1_Datao = 32'b0;
    reg signed [31:0] P1_P2_P1_EAX = 32'b0;
    reg signed [31:0] P1_P2_P1_EBX = 32'b0;
    reg P1_P2_P1_Extended = 1'b0;
    reg P1_P2_P1_Flush = 1'b0;
    reg P1_P2_P1_HOLD = 1'b0;
    reg signed [31:0] P1_P2_P1_InstAddrPointer = 32'b0;
    reg [7:0] P1_P2_P1_InstQueue [15:0];
    reg [4:0] P1_P2_P1_InstQueueRd_Addr = 5'b0;
    reg [4:0] P1_P2_P1_InstQueueWr_Addr = 5'b0;
    reg P1_P2_P1_M_IO_n = 1'b0;
    reg P1_P2_P1_MemoryFetch = 1'b0;
    reg P1_P2_P1_More = 1'b0;
    reg P1_P2_P1_NA_n = 1'b0;
    reg P1_P2_P1_NonAligned = 1'b0;
    reg signed [31:0] P1_P2_P1_PhyAddrPointer = 32'b0;
    reg P1_P2_P1_READY_n = 1'b0;
    reg P1_P2_P1_RESET = 1'b0;
    reg P1_P2_P1_ReadRequest = 1'b0;
    reg P1_P2_P1_RequestPending = 1'b0;
    reg [2:0] P1_P2_P1_State = 3'b0;
    reg [3:0] P1_P2_P1_State2 = 4'b0;
    reg P1_P2_P1_StateBS16 = 1'b0;
    reg P1_P2_P1_StateNA = 1'b0;
    reg P1_P2_P1_W_R_n = 1'b0;
    reg signed [31:0] P1_P2_P1_fWord = 32'b0;
    reg [15:0] P1_P2_P1_lWord = 16'b0;
    reg signed [31:0] P1_P2_P1_rEIP = 32'b0;
    reg [14:0] P1_P2_P1_uWord = 15'b0;
    reg P1_P2_P2_ADS_n = 1'b0;
    reg [29:0] P1_P2_P2_Address = 30'b0;
    reg [3:0] P1_P2_P2_BE_n = 4'b0;
    reg P1_P2_P2_BS16_n = 1'b0;
    reg [3:0] P1_P2_P2_ByteEnable = 4'b0;
    reg P1_P2_P2_CLOCK = 1'b0;
    reg P1_P2_P2_CodeFetch = 1'b0;
    reg P1_P2_P2_D_C_n = 1'b0;
    reg signed [31:0] P1_P2_P2_DataWidth = 32'b0;
    reg [31:0] P1_P2_P2_Datai = 32'b0;
    reg signed [31:0] P1_P2_P2_Datao = 32'b0;
    reg signed [31:0] P1_P2_P2_EAX = 32'b0;
    reg signed [31:0] P1_P2_P2_EBX = 32'b0;
    reg P1_P2_P2_Extended = 1'b0;
    reg P1_P2_P2_Flush = 1'b0;
    reg P1_P2_P2_HOLD = 1'b0;
    reg signed [31:0] P1_P2_P2_InstAddrPointer = 32'b0;
    reg [7:0] P1_P2_P2_InstQueue [15:0];
    reg [4:0] P1_P2_P2_InstQueueRd_Addr = 5'b0;
    reg [4:0] P1_P2_P2_InstQueueWr_Addr = 5'b0;
    reg P1_P2_P2_M_IO_n = 1'b0;
    reg P1_P2_P2_MemoryFetch = 1'b0;
    reg P1_P2_P2_More = 1'b0;
    reg P1_P2_P2_NA_n = 1'b0;
    reg P1_P2_P2_NonAligned = 1'b0;
    reg signed [31:0] P1_P2_P2_PhyAddrPointer = 32'b0;
    reg P1_P2_P2_READY_n = 1'b0;
    reg P1_P2_P2_RESET = 1'b0;
    reg P1_P2_P2_ReadRequest = 1'b0;
    reg P1_P2_P2_RequestPending = 1'b0;
    reg [2:0] P1_P2_P2_State = 3'b0;
    reg [3:0] P1_P2_P2_State2 = 4'b0;
    reg P1_P2_P2_StateBS16 = 1'b0;
    reg P1_P2_P2_StateNA = 1'b0;
    reg P1_P2_P2_W_R_n = 1'b0;
    reg signed [31:0] P1_P2_P2_fWord = 32'b0;
    reg [15:0] P1_P2_P2_lWord = 16'b0;
    reg signed [31:0] P1_P2_P2_rEIP = 32'b0;
    reg [14:0] P1_P2_P2_uWord = 15'b0;
    reg P1_P2_P3_ADS_n = 1'b0;
    reg [29:0] P1_P2_P3_Address = 30'b0;
    reg [3:0] P1_P2_P3_BE_n = 4'b0;
    reg P1_P2_P3_BS16_n = 1'b0;
    reg [3:0] P1_P2_P3_ByteEnable = 4'b0;
    reg P1_P2_P3_CLOCK = 1'b0;
    reg P1_P2_P3_CodeFetch = 1'b0;
    reg P1_P2_P3_D_C_n = 1'b0;
    reg signed [31:0] P1_P2_P3_DataWidth = 32'b0;
    reg [31:0] P1_P2_P3_Datai = 32'b0;
    reg signed [31:0] P1_P2_P3_Datao = 32'b0;
    reg signed [31:0] P1_P2_P3_EAX = 32'b0;
    reg signed [31:0] P1_P2_P3_EBX = 32'b0;
    reg P1_P2_P3_Extended = 1'b0;
    reg P1_P2_P3_Flush = 1'b0;
    reg P1_P2_P3_HOLD = 1'b0;
    reg signed [31:0] P1_P2_P3_InstAddrPointer = 32'b0;
    reg [7:0] P1_P2_P3_InstQueue [15:0];
    reg [4:0] P1_P2_P3_InstQueueRd_Addr = 5'b0;
    reg [4:0] P1_P2_P3_InstQueueWr_Addr = 5'b0;
    reg P1_P2_P3_M_IO_n = 1'b0;
    reg P1_P2_P3_MemoryFetch = 1'b0;
    reg P1_P2_P3_More = 1'b0;
    reg P1_P2_P3_NA_n = 1'b0;
    reg P1_P2_P3_NonAligned = 1'b0;
    reg signed [31:0] P1_P2_P3_PhyAddrPointer = 32'b0;
    reg P1_P2_P3_READY_n = 1'b0;
    reg P1_P2_P3_RESET = 1'b0;
    reg P1_P2_P3_ReadRequest = 1'b0;
    reg P1_P2_P3_RequestPending = 1'b0;
    reg [2:0] P1_P2_P3_State = 3'b0;
    reg [3:0] P1_P2_P3_State2 = 4'b0;
    reg P1_P2_P3_StateBS16 = 1'b0;
    reg P1_P2_P3_StateNA = 1'b0;
    reg P1_P2_P3_W_R_n = 1'b0;
    reg signed [31:0] P1_P2_P3_fWord = 32'b0;
    reg [15:0] P1_P2_P3_lWord = 16'b0;
    reg signed [31:0] P1_P2_P3_rEIP = 32'b0;
    reg [14:0] P1_P2_P3_uWord = 15'b0;
    reg [29:0] P1_P2_addr1 = 30'b0;
    reg [29:0] P1_P2_addr2 = 30'b0;
    reg [29:0] P1_P2_addr3 = 30'b0;
    reg [29:0] P1_P2_address1 = 30'b0;
    reg [29:0] P1_P2_address2 = 30'b0;
    reg P1_P2_ads1 = 1'b0;
    reg P1_P2_ads2 = 1'b0;
    reg P1_P2_ads3 = 1'b0;
    reg P1_P2_ast1 = 1'b0;
    reg P1_P2_ast2 = 1'b0;
    reg [3:0] P1_P2_be1 = 4'b0;
    reg [3:0] P1_P2_be2 = 4'b0;
    reg [3:0] P1_P2_be3 = 4'b0;
    reg P1_P2_bs16 = 1'b0;
    reg signed [31:0] P1_P2_buf1 = 32'b0;
    reg signed [31:0] P1_P2_buf2 = 32'b0;
    reg P1_P2_clock = 1'b0;
    reg [31:0] P1_P2_datai = 32'b0;
    reg signed [31:0] P1_P2_datao = 32'b0;
    reg P1_P2_dc = 1'b0;
    reg P1_P2_dc1 = 1'b0;
    reg P1_P2_dc2 = 1'b0;
    reg P1_P2_dc3 = 1'b0;
    reg signed [31:0] P1_P2_di1 = 32'b0;
    reg signed [31:0] P1_P2_di2 = 32'b0;
    reg signed [31:0] P1_P2_di3 = 32'b0;
    reg [31:0] P1_P2_do1 = 32'b0;
    reg [31:0] P1_P2_do2 = 32'b0;
    reg [31:0] P1_P2_do3 = 32'b0;
    reg P1_P2_hold = 1'b0;
    reg P1_P2_mio = 1'b0;
    reg P1_P2_mio1 = 1'b0;
    reg P1_P2_mio2 = 1'b0;
    reg P1_P2_mio3 = 1'b0;
    reg P1_P2_na = 1'b0;
    reg P1_P2_rdy1 = 1'b0;
    reg P1_P2_rdy2 = 1'b0;
    reg P1_P2_rdy3 = 1'b0;
    reg P1_P2_ready1 = 1'b0;
    reg P1_P2_ready11 = 1'b0;
    reg P1_P2_ready12 = 1'b0;
    reg P1_P2_ready2 = 1'b0;
    reg P1_P2_ready21 = 1'b0;
    reg P1_P2_ready22 = 1'b0;
    reg P1_P2_reset = 1'b0;
    reg P1_P2_wr = 1'b0;
    reg P1_P2_wr1 = 1'b0;
    reg P1_P2_wr2 = 1'b0;
    reg P1_P2_wr3 = 1'b0;
    reg P1_P3_B = 1'b0;
    reg signed [31:0] P1_P3_IR = 32'b0;
    reg [19:0] P1_P3_MAR = 20'b0;
    reg signed [31:0] P1_P3_MBR = 32'b0;
    reg [19:0] P1_P3_addr = 20'b0;
    reg P1_P3_cf = 1'b0;
    reg P1_P3_clock = 1'b0;
    reg signed [31:0] P1_P3_d = 32'b0;
    reg [31:0] P1_P3_datai = 32'b0;
    reg signed [31:0] P1_P3_datao = 32'b0;
    reg [2:0] P1_P3_df = 3'b0;
    reg [3:0] P1_P3_ff = 4'b0;
    reg signed [31:0] P1_P3_m = 32'b0;
    reg [1:0] P1_P3_mf = 2'b0;
    reg signed [31:0] P1_P3_r = 32'b0;
    reg P1_P3_rd = 1'b0;
    reg signed [31:0] P1_P3_reg0 = 32'b0;
    reg signed [31:0] P1_P3_reg1 = 32'b0;
    reg signed [31:0] P1_P3_reg2 = 32'b0;
    reg signed [31:0] P1_P3_reg3 = 32'b0;
    reg P1_P3_reset = 1'b0;
    reg [1:0] P1_P3_s = 2'b0;
    reg P1_P3_state = 1'b0;
    reg signed [31:0] P1_P3_t = 32'b0;
    reg [19:0] P1_P3_tail = 20'b0;
    reg signed [31:0] P1_P3_temp = 32'b0;
    reg P1_P3_wr = 1'b0;
    reg P1_P4_B = 1'b0;
    reg signed [31:0] P1_P4_IR = 32'b0;
    reg [19:0] P1_P4_MAR = 20'b0;
    reg signed [31:0] P1_P4_MBR = 32'b0;
    reg [19:0] P1_P4_addr = 20'b0;
    reg P1_P4_cf = 1'b0;
    reg P1_P4_clock = 1'b0;
    reg signed [31:0] P1_P4_d = 32'b0;
    reg [31:0] P1_P4_datai = 32'b0;
    reg signed [31:0] P1_P4_datao = 32'b0;
    reg [2:0] P1_P4_df = 3'b0;
    reg [3:0] P1_P4_ff = 4'b0;
    reg signed [31:0] P1_P4_m = 32'b0;
    reg [1:0] P1_P4_mf = 2'b0;
    reg signed [31:0] P1_P4_r = 32'b0;
    reg P1_P4_rd = 1'b0;
    reg signed [31:0] P1_P4_reg0 = 32'b0;
    reg signed [31:0] P1_P4_reg1 = 32'b0;
    reg signed [31:0] P1_P4_reg2 = 32'b0;
    reg signed [31:0] P1_P4_reg3 = 32'b0;
    reg P1_P4_reset = 1'b0;
    reg [1:0] P1_P4_s = 2'b0;
    reg P1_P4_state = 1'b0;
    reg signed [31:0] P1_P4_t = 32'b0;
    reg [19:0] P1_P4_tail = 20'b0;
    reg signed [31:0] P1_P4_temp = 32'b0;
    reg P1_P4_wr = 1'b0;
    reg [29:0] P1_ad11 = 30'b0;
    reg [29:0] P1_ad12 = 30'b0;
    reg [29:0] P1_ad21 = 30'b0;
    reg [29:0] P1_ad22 = 30'b0;
    reg [19:0] P1_ad31 = 20'b0;
    reg [19:0] P1_ad41 = 20'b0;
    reg P1_as11 = 1'b0;
    reg P1_as12 = 1'b0;
    reg P1_as21 = 1'b0;
    reg P1_as22 = 1'b0;
    reg [2:0] P1_aux = 3'b0;
    reg P1_bs = 1'b0;
    reg P1_clock = 1'b0;
    reg P1_dc1 = 1'b0;
    reg P1_dc2 = 1'b0;
    reg signed [31:0] P1_di1 = 32'b0;
    reg signed [31:0] P1_di2 = 32'b0;
    reg signed [31:0] P1_di3 = 32'b0;
    reg signed [31:0] P1_di4 = 32'b0;
    reg [31:0] P1_din = 32'b0;
    reg [31:0] P1_do1 = 32'b0;
    reg [31:0] P1_do2 = 32'b0;
    reg [31:0] P1_do3 = 32'b0;
    reg [31:0] P1_do4 = 32'b0;
    reg [19:0] P1_dout = 20'b0;
    reg P1_hold = 1'b0;
    reg P1_mio1 = 1'b0;
    reg P1_mio2 = 1'b0;
    reg P1_na = 1'b0;
    reg P1_r11 = 1'b0;
    reg P1_r12 = 1'b0;
    reg P1_r21 = 1'b0;
    reg P1_r22 = 1'b0;
    reg P1_rd3 = 1'b0;
    reg P1_rd4 = 1'b0;
    reg P1_reset = 1'b0;
    reg P1_sel = 1'b0;
    reg [29:0] P1_tad1 = 30'b0;
    reg [29:0] P1_tad2 = 30'b0;
    reg [19:0] P1_tad3 = 20'b0;
    reg [19:0] P1_tad4 = 20'b0;
    reg signed [31:0] P1_td1 = 32'b0;
    reg signed [31:0] P1_td2 = 32'b0;
    reg P1_wr1 = 1'b0;
    reg P1_wr2 = 1'b0;
    reg P1_wr3 = 1'b0;
    reg P1_wr4 = 1'b0;
    reg P2_P1_P1_ADS_n = 1'b0;
    reg [29:0] P2_P1_P1_Address = 30'b0;
    reg [3:0] P2_P1_P1_BE_n = 4'b0;
    reg P2_P1_P1_BS16_n = 1'b0;
    reg [3:0] P2_P1_P1_ByteEnable = 4'b0;
    reg P2_P1_P1_CLOCK = 1'b0;
    reg P2_P1_P1_CodeFetch = 1'b0;
    reg P2_P1_P1_D_C_n = 1'b0;
    reg signed [31:0] P2_P1_P1_DataWidth = 32'b0;
    reg [31:0] P2_P1_P1_Datai = 32'b0;
    reg signed [31:0] P2_P1_P1_Datao = 32'b0;
    reg signed [31:0] P2_P1_P1_EAX = 32'b0;
    reg signed [31:0] P2_P1_P1_EBX = 32'b0;
    reg P2_P1_P1_Extended = 1'b0;
    reg P2_P1_P1_Flush = 1'b0;
    reg P2_P1_P1_HOLD = 1'b0;
    reg signed [31:0] P2_P1_P1_InstAddrPointer = 32'b0;
    reg [7:0] P2_P1_P1_InstQueue [15:0];
    reg [4:0] P2_P1_P1_InstQueueRd_Addr = 5'b0;
    reg [4:0] P2_P1_P1_InstQueueWr_Addr = 5'b0;
    reg P2_P1_P1_M_IO_n = 1'b0;
    reg P2_P1_P1_MemoryFetch = 1'b0;
    reg P2_P1_P1_More = 1'b0;
    reg P2_P1_P1_NA_n = 1'b0;
    reg P2_P1_P1_NonAligned = 1'b0;
    reg signed [31:0] P2_P1_P1_PhyAddrPointer = 32'b0;
    reg P2_P1_P1_READY_n = 1'b0;
    reg P2_P1_P1_RESET = 1'b0;
    reg P2_P1_P1_ReadRequest = 1'b0;
    reg P2_P1_P1_RequestPending = 1'b0;
    reg [2:0] P2_P1_P1_State = 3'b0;
    reg [3:0] P2_P1_P1_State2 = 4'b0;
    reg P2_P1_P1_StateBS16 = 1'b0;
    reg P2_P1_P1_StateNA = 1'b0;
    reg P2_P1_P1_W_R_n = 1'b0;
    reg signed [31:0] P2_P1_P1_fWord = 32'b0;
    reg [15:0] P2_P1_P1_lWord = 16'b0;
    reg signed [31:0] P2_P1_P1_rEIP = 32'b0;
    reg [14:0] P2_P1_P1_uWord = 15'b0;
    reg P2_P1_P2_ADS_n = 1'b0;
    reg [29:0] P2_P1_P2_Address = 30'b0;
    reg [3:0] P2_P1_P2_BE_n = 4'b0;
    reg P2_P1_P2_BS16_n = 1'b0;
    reg [3:0] P2_P1_P2_ByteEnable = 4'b0;
    reg P2_P1_P2_CLOCK = 1'b0;
    reg P2_P1_P2_CodeFetch = 1'b0;
    reg P2_P1_P2_D_C_n = 1'b0;
    reg signed [31:0] P2_P1_P2_DataWidth = 32'b0;
    reg [31:0] P2_P1_P2_Datai = 32'b0;
    reg signed [31:0] P2_P1_P2_Datao = 32'b0;
    reg signed [31:0] P2_P1_P2_EAX = 32'b0;
    reg signed [31:0] P2_P1_P2_EBX = 32'b0;
    reg P2_P1_P2_Extended = 1'b0;
    reg P2_P1_P2_Flush = 1'b0;
    reg P2_P1_P2_HOLD = 1'b0;
    reg signed [31:0] P2_P1_P2_InstAddrPointer = 32'b0;
    reg [7:0] P2_P1_P2_InstQueue [15:0];
    reg [4:0] P2_P1_P2_InstQueueRd_Addr = 5'b0;
    reg [4:0] P2_P1_P2_InstQueueWr_Addr = 5'b0;
    reg P2_P1_P2_M_IO_n = 1'b0;
    reg P2_P1_P2_MemoryFetch = 1'b0;
    reg P2_P1_P2_More = 1'b0;
    reg P2_P1_P2_NA_n = 1'b0;
    reg P2_P1_P2_NonAligned = 1'b0;
    reg signed [31:0] P2_P1_P2_PhyAddrPointer = 32'b0;
    reg P2_P1_P2_READY_n = 1'b0;
    reg P2_P1_P2_RESET = 1'b0;
    reg P2_P1_P2_ReadRequest = 1'b0;
    reg P2_P1_P2_RequestPending = 1'b0;
    reg [2:0] P2_P1_P2_State = 3'b0;
    reg [3:0] P2_P1_P2_State2 = 4'b0;
    reg P2_P1_P2_StateBS16 = 1'b0;
    reg P2_P1_P2_StateNA = 1'b0;
    reg P2_P1_P2_W_R_n = 1'b0;
    reg signed [31:0] P2_P1_P2_fWord = 32'b0;
    reg [15:0] P2_P1_P2_lWord = 16'b0;
    reg signed [31:0] P2_P1_P2_rEIP = 32'b0;
    reg [14:0] P2_P1_P2_uWord = 15'b0;
    reg P2_P1_P3_ADS_n = 1'b0;
    reg [29:0] P2_P1_P3_Address = 30'b0;
    reg [3:0] P2_P1_P3_BE_n = 4'b0;
    reg P2_P1_P3_BS16_n = 1'b0;
    reg [3:0] P2_P1_P3_ByteEnable = 4'b0;
    reg P2_P1_P3_CLOCK = 1'b0;
    reg P2_P1_P3_CodeFetch = 1'b0;
    reg P2_P1_P3_D_C_n = 1'b0;
    reg signed [31:0] P2_P1_P3_DataWidth = 32'b0;
    reg [31:0] P2_P1_P3_Datai = 32'b0;
    reg signed [31:0] P2_P1_P3_Datao = 32'b0;
    reg signed [31:0] P2_P1_P3_EAX = 32'b0;
    reg signed [31:0] P2_P1_P3_EBX = 32'b0;
    reg P2_P1_P3_Extended = 1'b0;
    reg P2_P1_P3_Flush = 1'b0;
    reg P2_P1_P3_HOLD = 1'b0;
    reg signed [31:0] P2_P1_P3_InstAddrPointer = 32'b0;
    reg [7:0] P2_P1_P3_InstQueue [15:0];
    reg [4:0] P2_P1_P3_InstQueueRd_Addr = 5'b0;
    reg [4:0] P2_P1_P3_InstQueueWr_Addr = 5'b0;
    reg P2_P1_P3_M_IO_n = 1'b0;
    reg P2_P1_P3_MemoryFetch = 1'b0;
    reg P2_P1_P3_More = 1'b0;
    reg P2_P1_P3_NA_n = 1'b0;
    reg P2_P1_P3_NonAligned = 1'b0;
    reg signed [31:0] P2_P1_P3_PhyAddrPointer = 32'b0;
    reg P2_P1_P3_READY_n = 1'b0;
    reg P2_P1_P3_RESET = 1'b0;
    reg P2_P1_P3_ReadRequest = 1'b0;
    reg P2_P1_P3_RequestPending = 1'b0;
    reg [2:0] P2_P1_P3_State = 3'b0;
    reg [3:0] P2_P1_P3_State2 = 4'b0;
    reg P2_P1_P3_StateBS16 = 1'b0;
    reg P2_P1_P3_StateNA = 1'b0;
    reg P2_P1_P3_W_R_n = 1'b0;
    reg signed [31:0] P2_P1_P3_fWord = 32'b0;
    reg [15:0] P2_P1_P3_lWord = 16'b0;
    reg signed [31:0] P2_P1_P3_rEIP = 32'b0;
    reg [14:0] P2_P1_P3_uWord = 15'b0;
    reg [29:0] P2_P1_addr1 = 30'b0;
    reg [29:0] P2_P1_addr2 = 30'b0;
    reg [29:0] P2_P1_addr3 = 30'b0;
    reg [29:0] P2_P1_address1 = 30'b0;
    reg [29:0] P2_P1_address2 = 30'b0;
    reg P2_P1_ads1 = 1'b0;
    reg P2_P1_ads2 = 1'b0;
    reg P2_P1_ads3 = 1'b0;
    reg P2_P1_ast1 = 1'b0;
    reg P2_P1_ast2 = 1'b0;
    reg [3:0] P2_P1_be1 = 4'b0;
    reg [3:0] P2_P1_be2 = 4'b0;
    reg [3:0] P2_P1_be3 = 4'b0;
    reg P2_P1_bs16 = 1'b0;
    reg signed [31:0] P2_P1_buf1 = 32'b0;
    reg signed [31:0] P2_P1_buf2 = 32'b0;
    reg P2_P1_clock = 1'b0;
    reg [31:0] P2_P1_datai = 32'b0;
    reg signed [31:0] P2_P1_datao = 32'b0;
    reg P2_P1_dc = 1'b0;
    reg P2_P1_dc1 = 1'b0;
    reg P2_P1_dc2 = 1'b0;
    reg P2_P1_dc3 = 1'b0;
    reg signed [31:0] P2_P1_di1 = 32'b0;
    reg signed [31:0] P2_P1_di2 = 32'b0;
    reg signed [31:0] P2_P1_di3 = 32'b0;
    reg [31:0] P2_P1_do1 = 32'b0;
    reg [31:0] P2_P1_do2 = 32'b0;
    reg [31:0] P2_P1_do3 = 32'b0;
    reg P2_P1_hold = 1'b0;
    reg P2_P1_mio = 1'b0;
    reg P2_P1_mio1 = 1'b0;
    reg P2_P1_mio2 = 1'b0;
    reg P2_P1_mio3 = 1'b0;
    reg P2_P1_na = 1'b0;
    reg P2_P1_rdy1 = 1'b0;
    reg P2_P1_rdy2 = 1'b0;
    reg P2_P1_rdy3 = 1'b0;
    reg P2_P1_ready1 = 1'b0;
    reg P2_P1_ready11 = 1'b0;
    reg P2_P1_ready12 = 1'b0;
    reg P2_P1_ready2 = 1'b0;
    reg P2_P1_ready21 = 1'b0;
    reg P2_P1_ready22 = 1'b0;
    reg P2_P1_reset = 1'b0;
    reg P2_P1_wr = 1'b0;
    reg P2_P1_wr1 = 1'b0;
    reg P2_P1_wr2 = 1'b0;
    reg P2_P1_wr3 = 1'b0;
    reg P2_P2_P1_ADS_n = 1'b0;
    reg [29:0] P2_P2_P1_Address = 30'b0;
    reg [3:0] P2_P2_P1_BE_n = 4'b0;
    reg P2_P2_P1_BS16_n = 1'b0;
    reg [3:0] P2_P2_P1_ByteEnable = 4'b0;
    reg P2_P2_P1_CLOCK = 1'b0;
    reg P2_P2_P1_CodeFetch = 1'b0;
    reg P2_P2_P1_D_C_n = 1'b0;
    reg signed [31:0] P2_P2_P1_DataWidth = 32'b0;
    reg [31:0] P2_P2_P1_Datai = 32'b0;
    reg signed [31:0] P2_P2_P1_Datao = 32'b0;
    reg signed [31:0] P2_P2_P1_EAX = 32'b0;
    reg signed [31:0] P2_P2_P1_EBX = 32'b0;
    reg P2_P2_P1_Extended = 1'b0;
    reg P2_P2_P1_Flush = 1'b0;
    reg P2_P2_P1_HOLD = 1'b0;
    reg signed [31:0] P2_P2_P1_InstAddrPointer = 32'b0;
    reg [7:0] P2_P2_P1_InstQueue [15:0];
    reg [4:0] P2_P2_P1_InstQueueRd_Addr = 5'b0;
    reg [4:0] P2_P2_P1_InstQueueWr_Addr = 5'b0;
    reg P2_P2_P1_M_IO_n = 1'b0;
    reg P2_P2_P1_MemoryFetch = 1'b0;
    reg P2_P2_P1_More = 1'b0;
    reg P2_P2_P1_NA_n = 1'b0;
    reg P2_P2_P1_NonAligned = 1'b0;
    reg signed [31:0] P2_P2_P1_PhyAddrPointer = 32'b0;
    reg P2_P2_P1_READY_n = 1'b0;
    reg P2_P2_P1_RESET = 1'b0;
    reg P2_P2_P1_ReadRequest = 1'b0;
    reg P2_P2_P1_RequestPending = 1'b0;
    reg [2:0] P2_P2_P1_State = 3'b0;
    reg [3:0] P2_P2_P1_State2 = 4'b0;
    reg P2_P2_P1_StateBS16 = 1'b0;
    reg P2_P2_P1_StateNA = 1'b0;
    reg P2_P2_P1_W_R_n = 1'b0;
    reg signed [31:0] P2_P2_P1_fWord = 32'b0;
    reg [15:0] P2_P2_P1_lWord = 16'b0;
    reg signed [31:0] P2_P2_P1_rEIP = 32'b0;
    reg [14:0] P2_P2_P1_uWord = 15'b0;
    reg P2_P2_P2_ADS_n = 1'b0;
    reg [29:0] P2_P2_P2_Address = 30'b0;
    reg [3:0] P2_P2_P2_BE_n = 4'b0;
    reg P2_P2_P2_BS16_n = 1'b0;
    reg [3:0] P2_P2_P2_ByteEnable = 4'b0;
    reg P2_P2_P2_CLOCK = 1'b0;
    reg P2_P2_P2_CodeFetch = 1'b0;
    reg P2_P2_P2_D_C_n = 1'b0;
    reg signed [31:0] P2_P2_P2_DataWidth = 32'b0;
    reg [31:0] P2_P2_P2_Datai = 32'b0;
    reg signed [31:0] P2_P2_P2_Datao = 32'b0;
    reg signed [31:0] P2_P2_P2_EAX = 32'b0;
    reg signed [31:0] P2_P2_P2_EBX = 32'b0;
    reg P2_P2_P2_Extended = 1'b0;
    reg P2_P2_P2_Flush = 1'b0;
    reg P2_P2_P2_HOLD = 1'b0;
    reg signed [31:0] P2_P2_P2_InstAddrPointer = 32'b0;
    reg [7:0] P2_P2_P2_InstQueue [15:0];
    reg [4:0] P2_P2_P2_InstQueueRd_Addr = 5'b0;
    reg [4:0] P2_P2_P2_InstQueueWr_Addr = 5'b0;
    reg P2_P2_P2_M_IO_n = 1'b0;
    reg P2_P2_P2_MemoryFetch = 1'b0;
    reg P2_P2_P2_More = 1'b0;
    reg P2_P2_P2_NA_n = 1'b0;
    reg P2_P2_P2_NonAligned = 1'b0;
    reg signed [31:0] P2_P2_P2_PhyAddrPointer = 32'b0;
    reg P2_P2_P2_READY_n = 1'b0;
    reg P2_P2_P2_RESET = 1'b0;
    reg P2_P2_P2_ReadRequest = 1'b0;
    reg P2_P2_P2_RequestPending = 1'b0;
    reg [2:0] P2_P2_P2_State = 3'b0;
    reg [3:0] P2_P2_P2_State2 = 4'b0;
    reg P2_P2_P2_StateBS16 = 1'b0;
    reg P2_P2_P2_StateNA = 1'b0;
    reg P2_P2_P2_W_R_n = 1'b0;
    reg signed [31:0] P2_P2_P2_fWord = 32'b0;
    reg [15:0] P2_P2_P2_lWord = 16'b0;
    reg signed [31:0] P2_P2_P2_rEIP = 32'b0;
    reg [14:0] P2_P2_P2_uWord = 15'b0;
    reg P2_P2_P3_ADS_n = 1'b0;
    reg [29:0] P2_P2_P3_Address = 30'b0;
    reg [3:0] P2_P2_P3_BE_n = 4'b0;
    reg P2_P2_P3_BS16_n = 1'b0;
    reg [3:0] P2_P2_P3_ByteEnable = 4'b0;
    reg P2_P2_P3_CLOCK = 1'b0;
    reg P2_P2_P3_CodeFetch = 1'b0;
    reg P2_P2_P3_D_C_n = 1'b0;
    reg signed [31:0] P2_P2_P3_DataWidth = 32'b0;
    reg [31:0] P2_P2_P3_Datai = 32'b0;
    reg signed [31:0] P2_P2_P3_Datao = 32'b0;
    reg signed [31:0] P2_P2_P3_EAX = 32'b0;
    reg signed [31:0] P2_P2_P3_EBX = 32'b0;
    reg P2_P2_P3_Extended = 1'b0;
    reg P2_P2_P3_Flush = 1'b0;
    reg P2_P2_P3_HOLD = 1'b0;
    reg signed [31:0] P2_P2_P3_InstAddrPointer = 32'b0;
    reg [7:0] P2_P2_P3_InstQueue [15:0];
    reg [4:0] P2_P2_P3_InstQueueRd_Addr = 5'b0;
    reg [4:0] P2_P2_P3_InstQueueWr_Addr = 5'b0;
    reg P2_P2_P3_M_IO_n = 1'b0;
    reg P2_P2_P3_MemoryFetch = 1'b0;
    reg P2_P2_P3_More = 1'b0;
    reg P2_P2_P3_NA_n = 1'b0;
    reg P2_P2_P3_NonAligned = 1'b0;
    reg signed [31:0] P2_P2_P3_PhyAddrPointer = 32'b0;
    reg P2_P2_P3_READY_n = 1'b0;
    reg P2_P2_P3_RESET = 1'b0;
    reg P2_P2_P3_ReadRequest = 1'b0;
    reg P2_P2_P3_RequestPending = 1'b0;
    reg [2:0] P2_P2_P3_State = 3'b0;
    reg [3:0] P2_P2_P3_State2 = 4'b0;
    reg P2_P2_P3_StateBS16 = 1'b0;
    reg P2_P2_P3_StateNA = 1'b0;
    reg P2_P2_P3_W_R_n = 1'b0;
    reg signed [31:0] P2_P2_P3_fWord = 32'b0;
    reg [15:0] P2_P2_P3_lWord = 16'b0;
    reg signed [31:0] P2_P2_P3_rEIP = 32'b0;
    reg [14:0] P2_P2_P3_uWord = 15'b0;
    reg [29:0] P2_P2_addr1 = 30'b0;
    reg [29:0] P2_P2_addr2 = 30'b0;
    reg [29:0] P2_P2_addr3 = 30'b0;
    reg [29:0] P2_P2_address1 = 30'b0;
    reg [29:0] P2_P2_address2 = 30'b0;
    reg P2_P2_ads1 = 1'b0;
    reg P2_P2_ads2 = 1'b0;
    reg P2_P2_ads3 = 1'b0;
    reg P2_P2_ast1 = 1'b0;
    reg P2_P2_ast2 = 1'b0;
    reg [3:0] P2_P2_be1 = 4'b0;
    reg [3:0] P2_P2_be2 = 4'b0;
    reg [3:0] P2_P2_be3 = 4'b0;
    reg P2_P2_bs16 = 1'b0;
    reg signed [31:0] P2_P2_buf1 = 32'b0;
    reg signed [31:0] P2_P2_buf2 = 32'b0;
    reg P2_P2_clock = 1'b0;
    reg [31:0] P2_P2_datai = 32'b0;
    reg signed [31:0] P2_P2_datao = 32'b0;
    reg P2_P2_dc = 1'b0;
    reg P2_P2_dc1 = 1'b0;
    reg P2_P2_dc2 = 1'b0;
    reg P2_P2_dc3 = 1'b0;
    reg signed [31:0] P2_P2_di1 = 32'b0;
    reg signed [31:0] P2_P2_di2 = 32'b0;
    reg signed [31:0] P2_P2_di3 = 32'b0;
    reg [31:0] P2_P2_do1 = 32'b0;
    reg [31:0] P2_P2_do2 = 32'b0;
    reg [31:0] P2_P2_do3 = 32'b0;
    reg P2_P2_hold = 1'b0;
    reg P2_P2_mio = 1'b0;
    reg P2_P2_mio1 = 1'b0;
    reg P2_P2_mio2 = 1'b0;
    reg P2_P2_mio3 = 1'b0;
    reg P2_P2_na = 1'b0;
    reg P2_P2_rdy1 = 1'b0;
    reg P2_P2_rdy2 = 1'b0;
    reg P2_P2_rdy3 = 1'b0;
    reg P2_P2_ready1 = 1'b0;
    reg P2_P2_ready11 = 1'b0;
    reg P2_P2_ready12 = 1'b0;
    reg P2_P2_ready2 = 1'b0;
    reg P2_P2_ready21 = 1'b0;
    reg P2_P2_ready22 = 1'b0;
    reg P2_P2_reset = 1'b0;
    reg P2_P2_wr = 1'b0;
    reg P2_P2_wr1 = 1'b0;
    reg P2_P2_wr2 = 1'b0;
    reg P2_P2_wr3 = 1'b0;
    reg P2_P3_B = 1'b0;
    reg signed [31:0] P2_P3_IR = 32'b0;
    reg [19:0] P2_P3_MAR = 20'b0;
    reg signed [31:0] P2_P3_MBR = 32'b0;
    reg [19:0] P2_P3_addr = 20'b0;
    reg P2_P3_cf = 1'b0;
    reg P2_P3_clock = 1'b0;
    reg signed [31:0] P2_P3_d = 32'b0;
    reg [31:0] P2_P3_datai = 32'b0;
    reg signed [31:0] P2_P3_datao = 32'b0;
    reg [2:0] P2_P3_df = 3'b0;
    reg [3:0] P2_P3_ff = 4'b0;
    reg signed [31:0] P2_P3_m = 32'b0;
    reg [1:0] P2_P3_mf = 2'b0;
    reg signed [31:0] P2_P3_r = 32'b0;
    reg P2_P3_rd = 1'b0;
    reg signed [31:0] P2_P3_reg0 = 32'b0;
    reg signed [31:0] P2_P3_reg1 = 32'b0;
    reg signed [31:0] P2_P3_reg2 = 32'b0;
    reg signed [31:0] P2_P3_reg3 = 32'b0;
    reg P2_P3_reset = 1'b0;
    reg [1:0] P2_P3_s = 2'b0;
    reg P2_P3_state = 1'b0;
    reg signed [31:0] P2_P3_t = 32'b0;
    reg [19:0] P2_P3_tail = 20'b0;
    reg signed [31:0] P2_P3_temp = 32'b0;
    reg P2_P3_wr = 1'b0;
    reg P2_P4_B = 1'b0;
    reg signed [31:0] P2_P4_IR = 32'b0;
    reg [19:0] P2_P4_MAR = 20'b0;
    reg signed [31:0] P2_P4_MBR = 32'b0;
    reg [19:0] P2_P4_addr = 20'b0;
    reg P2_P4_cf = 1'b0;
    reg P2_P4_clock = 1'b0;
    reg signed [31:0] P2_P4_d = 32'b0;
    reg [31:0] P2_P4_datai = 32'b0;
    reg signed [31:0] P2_P4_datao = 32'b0;
    reg [2:0] P2_P4_df = 3'b0;
    reg [3:0] P2_P4_ff = 4'b0;
    reg signed [31:0] P2_P4_m = 32'b0;
    reg [1:0] P2_P4_mf = 2'b0;
    reg signed [31:0] P2_P4_r = 32'b0;
    reg P2_P4_rd = 1'b0;
    reg signed [31:0] P2_P4_reg0 = 32'b0;
    reg signed [31:0] P2_P4_reg1 = 32'b0;
    reg signed [31:0] P2_P4_reg2 = 32'b0;
    reg signed [31:0] P2_P4_reg3 = 32'b0;
    reg P2_P4_reset = 1'b0;
    reg [1:0] P2_P4_s = 2'b0;
    reg P2_P4_state = 1'b0;
    reg signed [31:0] P2_P4_t = 32'b0;
    reg [19:0] P2_P4_tail = 20'b0;
    reg signed [31:0] P2_P4_temp = 32'b0;
    reg P2_P4_wr = 1'b0;
    reg [29:0] P2_ad11 = 30'b0;
    reg [29:0] P2_ad12 = 30'b0;
    reg [29:0] P2_ad21 = 30'b0;
    reg [29:0] P2_ad22 = 30'b0;
    reg [19:0] P2_ad31 = 20'b0;
    reg [19:0] P2_ad41 = 20'b0;
    reg P2_as11 = 1'b0;
    reg P2_as12 = 1'b0;
    reg P2_as21 = 1'b0;
    reg P2_as22 = 1'b0;
    reg [2:0] P2_aux = 3'b0;
    reg P2_bs = 1'b0;
    reg P2_clock = 1'b0;
    reg P2_dc1 = 1'b0;
    reg P2_dc2 = 1'b0;
    reg signed [31:0] P2_di1 = 32'b0;
    reg signed [31:0] P2_di2 = 32'b0;
    reg signed [31:0] P2_di3 = 32'b0;
    reg signed [31:0] P2_di4 = 32'b0;
    reg [31:0] P2_din = 32'b0;
    reg [31:0] P2_do1 = 32'b0;
    reg [31:0] P2_do2 = 32'b0;
    reg [31:0] P2_do3 = 32'b0;
    reg [31:0] P2_do4 = 32'b0;
    reg [19:0] P2_dout = 20'b0;
    reg P2_hold = 1'b0;
    reg P2_mio1 = 1'b0;
    reg P2_mio2 = 1'b0;
    reg P2_na = 1'b0;
    reg P2_r11 = 1'b0;
    reg P2_r12 = 1'b0;
    reg P2_r21 = 1'b0;
    reg P2_r22 = 1'b0;
    reg P2_rd3 = 1'b0;
    reg P2_rd4 = 1'b0;
    reg P2_reset = 1'b0;
    reg P2_sel = 1'b0;
    reg [29:0] P2_tad1 = 30'b0;
    reg [29:0] P2_tad2 = 30'b0;
    reg [19:0] P2_tad3 = 20'b0;
    reg [19:0] P2_tad4 = 20'b0;
    reg signed [31:0] P2_td1 = 32'b0;
    reg signed [31:0] P2_td2 = 32'b0;
    reg P2_wr1 = 1'b0;
    reg P2_wr2 = 1'b0;
    reg P2_wr3 = 1'b0;
    reg P2_wr4 = 1'b0;
    reg [2:0] ax1 = 3'b0;
    reg [2:0] ax2 = 3'b0;
    reg signed [31:0] di1 = 32'b0;
    reg signed [31:0] di2 = 32'b0;
    reg [19:0] do1 = 20'b0;
    reg [19:0] do2 = 20'b0;
    reg [29:0] ris = 30'b0;
    reg sel1 = 1'b0;
    reg sel2 = 1'b0;

    always @(*) begin
        P1_clock = clock; $display(";A 0");		//(= P1_clock    clock )) ;0
    end

    always @(*) begin
        P1_reset = reset;    end

    always @(*) begin
        P1_hold = hold; $display(";A 2");		//(= P1_hold    hold )) ;2
    end

    always @(*) begin
        P1_na = na; $display(";A 3");		//(= P1_na    na )) ;3
    end

    always @(*) begin
        P1_bs = bs; $display(";A 4");		//(= P1_bs    bs )) ;4
    end

    always @(*) begin
        P1_sel = sel1; $display(";A 5");		//(= P1_sel    sel1 )) ;5
    end

    always @(*) begin
        do1 = P1_dout; $display(";A 6");		//(= do1    P1_dout )) ;6
    end

    always @(*) begin
        P1_din = di1; $display(";A 7");		//(= P1_din    di1 )) ;7
    end

    always @(*) begin
        ax1 = P1_aux; $display(";A 8");		//(= ax1    P1_aux )) ;8
    end

    always @(*) begin
        P1_P1_clock = P1_clock; $display(";A 9");		//(= P1_P1_clock    P1_clock )) ;9
    end

    always @(*) begin
        P1_P1_reset = P1_reset;    end

    always @(*) begin
        P1_P1_datai = P1_di1; $display(";A 11");		//(= P1_P1_datai    P1_di1 )) ;11
    end

    always @(*) begin
        P1_do1 = P1_P1_datao; $display(";A 12");		//(= P1_do1    P1_P1_datao )) ;12
    end

    always @(*) begin
        P1_P1_hold = P1_hold; $display(";A 13");		//(= P1_P1_hold    P1_hold )) ;13
    end

    always @(*) begin
        P1_P1_na = P1_na; $display(";A 14");		//(= P1_P1_na    P1_na )) ;14
    end

    always @(*) begin
        P1_P1_bs16 = P1_bs; $display(";A 15");		//(= P1_P1_bs16    P1_bs )) ;15
    end

    always @(*) begin
        P1_ad11 = P1_P1_address1; $display(";A 16");		//(= P1_ad11    P1_P1_address1 )) ;16
    end

    always @(*) begin
        P1_ad12 = P1_P1_address2; $display(";A 17");		//(= P1_ad12    P1_P1_address2 )) ;17
    end

    always @(*) begin
        P1_wr1 = P1_P1_wr; $display(";A 18");		//(= P1_wr1    P1_P1_wr )) ;18
    end

    always @(*) begin
        P1_dc1 = P1_P1_dc; $display(";A 19");		//(= P1_dc1    P1_P1_dc )) ;19
    end

    always @(*) begin
        P1_mio1 = P1_P1_mio; $display(";A 20");		//(= P1_mio1    P1_P1_mio )) ;20
    end

    always @(*) begin
        P1_as11 = P1_P1_ast1; $display(";A 21");		//(= P1_as11    P1_P1_ast1 )) ;21
    end

    always @(*) begin
        P1_as12 = P1_P1_ast2; $display(";A 22");		//(= P1_as12    P1_P1_ast2 )) ;22
    end

    always @(*) begin
        P1_P1_ready1 = P1_r11; $display(";A 23");		//(= P1_P1_ready1    P1_r11 )) ;23
    end

    always @(*) begin
        P1_P1_ready2 = P1_r12; $display(";A 24");		//(= P1_P1_ready2    P1_r12 )) ;24
    end

    always @(*) begin
        P1_P1_be1 = P1_P1_P1_BE_n; $display(";A 25");		//(= P1_P1_be1    P1_P1_P1_BE_n )) ;25
    end

    always @(*) begin
        P1_P1_addr1 = P1_P1_P1_Address; $display(";A 26");		//(= P1_P1_addr1    P1_P1_P1_Address )) ;26
    end

    always @(*) begin
        P1_P1_wr1 = P1_P1_P1_W_R_n; $display(";A 27");		//(= P1_P1_wr1    P1_P1_P1_W_R_n )) ;27
    end

    always @(*) begin
        P1_P1_dc1 = P1_P1_P1_D_C_n; $display(";A 28");		//(= P1_P1_dc1    P1_P1_P1_D_C_n )) ;28
    end

    always @(*) begin
        P1_P1_mio1 = P1_P1_P1_M_IO_n; $display(";A 29");		//(= P1_P1_mio1    P1_P1_P1_M_IO_n )) ;29
    end

    always @(*) begin
        P1_P1_ads1 = P1_P1_P1_ADS_n; $display(";A 30");		//(= P1_P1_ads1    P1_P1_P1_ADS_n )) ;30
    end

    always @(*) begin
        P1_P1_P1_Datai = P1_P1_di1; $display(";A 31");		//(= P1_P1_P1_Datai    P1_P1_di1 )) ;31
    end

    always @(*) begin
        P1_P1_do1 = P1_P1_P1_Datao; $display(";A 32");		//(= P1_P1_do1    P1_P1_P1_Datao )) ;32
    end

    always @(*) begin
        P1_P1_P1_CLOCK = P1_P1_clock; $display(";A 33");		//(= P1_P1_P1_CLOCK    P1_P1_clock )) ;33
    end

    always @(*) begin
        P1_P1_P1_NA_n = P1_P1_na; $display(";A 34");		//(= P1_P1_P1_NA_n    P1_P1_na )) ;34
    end

    always @(*) begin
        P1_P1_P1_BS16_n = P1_P1_bs16; $display(";A 35");		//(= P1_P1_P1_BS16_n    P1_P1_bs16 )) ;35
    end

    always @(*) begin
        P1_P1_P1_READY_n = P1_P1_rdy1; $display(";A 36");		//(= P1_P1_P1_READY_n    P1_P1_rdy1 )) ;36
    end

    always @(*) begin
        P1_P1_P1_HOLD = P1_P1_hold; $display(";A 37");		//(= P1_P1_P1_HOLD    P1_P1_hold )) ;37
    end

    always @(*) begin
        P1_P1_P1_RESET = P1_P1_reset;    end

    always @(*) begin
        P1_P1_be2 = P1_P1_P2_BE_n; $display(";A 39");		//(= P1_P1_be2    P1_P1_P2_BE_n )) ;39
    end

    always @(*) begin
        P1_P1_addr2 = P1_P1_P2_Address; $display(";A 40");		//(= P1_P1_addr2    P1_P1_P2_Address )) ;40
    end

    always @(*) begin
        P1_P1_wr2 = P1_P1_P2_W_R_n; $display(";A 41");		//(= P1_P1_wr2    P1_P1_P2_W_R_n )) ;41
    end

    always @(*) begin
        P1_P1_dc2 = P1_P1_P2_D_C_n; $display(";A 42");		//(= P1_P1_dc2    P1_P1_P2_D_C_n )) ;42
    end

    always @(*) begin
        P1_P1_mio2 = P1_P1_P2_M_IO_n; $display(";A 43");		//(= P1_P1_mio2    P1_P1_P2_M_IO_n )) ;43
    end

    always @(*) begin
        P1_P1_ads2 = P1_P1_P2_ADS_n; $display(";A 44");		//(= P1_P1_ads2    P1_P1_P2_ADS_n )) ;44
    end

    always @(*) begin
        P1_P1_P2_Datai = P1_P1_di2; $display(";A 45");		//(= P1_P1_P2_Datai    P1_P1_di2 )) ;45
    end

    always @(*) begin
        P1_P1_do2 = P1_P1_P2_Datao; $display(";A 46");		//(= P1_P1_do2    P1_P1_P2_Datao )) ;46
    end

    always @(*) begin
        P1_P1_P2_CLOCK = P1_P1_clock; $display(";A 47");		//(= P1_P1_P2_CLOCK    P1_P1_clock )) ;47
    end

    always @(*) begin
        P1_P1_P2_NA_n = P1_P1_na; $display(";A 48");		//(= P1_P1_P2_NA_n    P1_P1_na )) ;48
    end

    always @(*) begin
        P1_P1_P2_BS16_n = P1_P1_bs16; $display(";A 49");		//(= P1_P1_P2_BS16_n    P1_P1_bs16 )) ;49
    end

    always @(*) begin
        P1_P1_P2_READY_n = P1_P1_rdy2; $display(";A 50");		//(= P1_P1_P2_READY_n    P1_P1_rdy2 )) ;50
    end

    always @(*) begin
        P1_P1_P2_HOLD = P1_P1_hold; $display(";A 51");		//(= P1_P1_P2_HOLD    P1_P1_hold )) ;51
    end

    always @(*) begin
        P1_P1_P2_RESET = P1_P1_reset;    end

    always @(*) begin
        P1_P1_be3 = P1_P1_P3_BE_n; $display(";A 53");		//(= P1_P1_be3    P1_P1_P3_BE_n )) ;53
    end

    always @(*) begin
        P1_P1_addr3 = P1_P1_P3_Address; $display(";A 54");		//(= P1_P1_addr3    P1_P1_P3_Address )) ;54
    end

    always @(*) begin
        P1_P1_wr3 = P1_P1_P3_W_R_n; $display(";A 55");		//(= P1_P1_wr3    P1_P1_P3_W_R_n )) ;55
    end

    always @(*) begin
        P1_P1_dc3 = P1_P1_P3_D_C_n; $display(";A 56");		//(= P1_P1_dc3    P1_P1_P3_D_C_n )) ;56
    end

    always @(*) begin
        P1_P1_mio3 = P1_P1_P3_M_IO_n; $display(";A 57");		//(= P1_P1_mio3    P1_P1_P3_M_IO_n )) ;57
    end

    always @(*) begin
        P1_P1_ads3 = P1_P1_P3_ADS_n; $display(";A 58");		//(= P1_P1_ads3    P1_P1_P3_ADS_n )) ;58
    end

    always @(*) begin
        P1_P1_P3_Datai = P1_P1_di3; $display(";A 59");		//(= P1_P1_P3_Datai    P1_P1_di3 )) ;59
    end

    always @(*) begin
        P1_P1_do3 = P1_P1_P3_Datao; $display(";A 60");		//(= P1_P1_do3    P1_P1_P3_Datao )) ;60
    end

    always @(*) begin
        P1_P1_P3_CLOCK = P1_P1_clock; $display(";A 61");		//(= P1_P1_P3_CLOCK    P1_P1_clock )) ;61
    end

    always @(*) begin
        P1_P1_P3_NA_n = P1_P1_na; $display(";A 62");		//(= P1_P1_P3_NA_n    P1_P1_na )) ;62
    end

    always @(*) begin
        P1_P1_P3_BS16_n = P1_P1_bs16; $display(";A 63");		//(= P1_P1_P3_BS16_n    P1_P1_bs16 )) ;63
    end

    always @(*) begin
        P1_P1_P3_READY_n = P1_P1_rdy3; $display(";A 64");		//(= P1_P1_P3_READY_n    P1_P1_rdy3 )) ;64
    end

    always @(*) begin
        P1_P1_P3_HOLD = P1_P1_hold; $display(";A 65");		//(= P1_P1_P3_HOLD    P1_P1_hold )) ;65
    end

    always @(*) begin
        P1_P1_P3_RESET = P1_P1_reset;    end

    always @(*) begin
        P1_P2_clock = P1_clock; $display(";A 67");		//(= P1_P2_clock    P1_clock )) ;67
    end

    always @(*) begin
        P1_P2_reset = P1_reset;    end

    always @(*) begin
        P1_P2_datai = P1_di2; $display(";A 69");		//(= P1_P2_datai    P1_di2 )) ;69
    end

    always @(*) begin
        P1_do2 = P1_P2_datao; $display(";A 70");		//(= P1_do2    P1_P2_datao )) ;70
    end

    always @(*) begin
        P1_P2_hold = P1_hold; $display(";A 71");		//(= P1_P2_hold    P1_hold )) ;71
    end

    always @(*) begin
        P1_P2_na = P1_na; $display(";A 72");		//(= P1_P2_na    P1_na )) ;72
    end

    always @(*) begin
        P1_P2_bs16 = P1_bs; $display(";A 73");		//(= P1_P2_bs16    P1_bs )) ;73
    end

    always @(*) begin
        P1_ad21 = P1_P2_address1; $display(";A 74");		//(= P1_ad21    P1_P2_address1 )) ;74
    end

    always @(*) begin
        P1_ad22 = P1_P2_address2; $display(";A 75");		//(= P1_ad22    P1_P2_address2 )) ;75
    end

    always @(*) begin
        P1_wr2 = P1_P2_wr; $display(";A 76");		//(= P1_wr2    P1_P2_wr )) ;76
    end

    always @(*) begin
        P1_dc2 = P1_P2_dc; $display(";A 77");		//(= P1_dc2    P1_P2_dc )) ;77
    end

    always @(*) begin
        P1_mio2 = P1_P2_mio; $display(";A 78");		//(= P1_mio2    P1_P2_mio )) ;78
    end

    always @(*) begin
        P1_as21 = P1_P2_ast1; $display(";A 79");		//(= P1_as21    P1_P2_ast1 )) ;79
    end

    always @(*) begin
        P1_as22 = P1_P2_ast2; $display(";A 80");		//(= P1_as22    P1_P2_ast2 )) ;80
    end

    always @(*) begin
        P1_P2_ready1 = P1_r21; $display(";A 81");		//(= P1_P2_ready1    P1_r21 )) ;81
    end

    always @(*) begin
        P1_P2_ready2 = P1_r22; $display(";A 82");		//(= P1_P2_ready2    P1_r22 )) ;82
    end

    always @(*) begin
        P1_P2_be1 = P1_P2_P1_BE_n; $display(";A 83");		//(= P1_P2_be1    P1_P2_P1_BE_n )) ;83
    end

    always @(*) begin
        P1_P2_addr1 = P1_P2_P1_Address; $display(";A 84");		//(= P1_P2_addr1    P1_P2_P1_Address )) ;84
    end

    always @(*) begin
        P1_P2_wr1 = P1_P2_P1_W_R_n; $display(";A 85");		//(= P1_P2_wr1    P1_P2_P1_W_R_n )) ;85
    end

    always @(*) begin
        P1_P2_dc1 = P1_P2_P1_D_C_n; $display(";A 86");		//(= P1_P2_dc1    P1_P2_P1_D_C_n )) ;86
    end

    always @(*) begin
        P1_P2_mio1 = P1_P2_P1_M_IO_n; $display(";A 87");		//(= P1_P2_mio1    P1_P2_P1_M_IO_n )) ;87
    end

    always @(*) begin
        P1_P2_ads1 = P1_P2_P1_ADS_n; $display(";A 88");		//(= P1_P2_ads1    P1_P2_P1_ADS_n )) ;88
    end

    always @(*) begin
        P1_P2_P1_Datai = P1_P2_di1; $display(";A 89");		//(= P1_P2_P1_Datai    P1_P2_di1 )) ;89
    end

    always @(*) begin
        P1_P2_do1 = P1_P2_P1_Datao; $display(";A 90");		//(= P1_P2_do1    P1_P2_P1_Datao )) ;90
    end

    always @(*) begin
        P1_P2_P1_CLOCK = P1_P2_clock; $display(";A 91");		//(= P1_P2_P1_CLOCK    P1_P2_clock )) ;91
    end

    always @(*) begin
        P1_P2_P1_NA_n = P1_P2_na; $display(";A 92");		//(= P1_P2_P1_NA_n    P1_P2_na )) ;92
    end

    always @(*) begin
        P1_P2_P1_BS16_n = P1_P2_bs16; $display(";A 93");		//(= P1_P2_P1_BS16_n    P1_P2_bs16 )) ;93
    end

    always @(*) begin
        P1_P2_P1_READY_n = P1_P2_rdy1; $display(";A 94");		//(= P1_P2_P1_READY_n    P1_P2_rdy1 )) ;94
    end

    always @(*) begin
        P1_P2_P1_HOLD = P1_P2_hold; $display(";A 95");		//(= P1_P2_P1_HOLD    P1_P2_hold )) ;95
    end

    always @(*) begin
        P1_P2_P1_RESET = P1_P2_reset;    end

    always @(*) begin
        P1_P2_be2 = P1_P2_P2_BE_n; $display(";A 97");		//(= P1_P2_be2    P1_P2_P2_BE_n )) ;97
    end

    always @(*) begin
        P1_P2_addr2 = P1_P2_P2_Address; $display(";A 98");		//(= P1_P2_addr2    P1_P2_P2_Address )) ;98
    end

    always @(*) begin
        P1_P2_wr2 = P1_P2_P2_W_R_n; $display(";A 99");		//(= P1_P2_wr2    P1_P2_P2_W_R_n )) ;99
    end

    always @(*) begin
        P1_P2_dc2 = P1_P2_P2_D_C_n; $display(";A 100");		//(= P1_P2_dc2    P1_P2_P2_D_C_n )) ;100
    end

    always @(*) begin
        P1_P2_mio2 = P1_P2_P2_M_IO_n; $display(";A 101");		//(= P1_P2_mio2    P1_P2_P2_M_IO_n )) ;101
    end

    always @(*) begin
        P1_P2_ads2 = P1_P2_P2_ADS_n; $display(";A 102");		//(= P1_P2_ads2    P1_P2_P2_ADS_n )) ;102
    end

    always @(*) begin
        P1_P2_P2_Datai = P1_P2_di2; $display(";A 103");		//(= P1_P2_P2_Datai    P1_P2_di2 )) ;103
    end

    always @(*) begin
        P1_P2_do2 = P1_P2_P2_Datao; $display(";A 104");		//(= P1_P2_do2    P1_P2_P2_Datao )) ;104
    end

    always @(*) begin
        P1_P2_P2_CLOCK = P1_P2_clock; $display(";A 105");		//(= P1_P2_P2_CLOCK    P1_P2_clock )) ;105
    end

    always @(*) begin
        P1_P2_P2_NA_n = P1_P2_na; $display(";A 106");		//(= P1_P2_P2_NA_n    P1_P2_na )) ;106
    end

    always @(*) begin
        P1_P2_P2_BS16_n = P1_P2_bs16; $display(";A 107");		//(= P1_P2_P2_BS16_n    P1_P2_bs16 )) ;107
    end

    always @(*) begin
        P1_P2_P2_READY_n = P1_P2_rdy2; $display(";A 108");		//(= P1_P2_P2_READY_n    P1_P2_rdy2 )) ;108
    end

    always @(*) begin
        P1_P2_P2_HOLD = P1_P2_hold; $display(";A 109");		//(= P1_P2_P2_HOLD    P1_P2_hold )) ;109
    end

    always @(*) begin
        P1_P2_P2_RESET = P1_P2_reset;    end

    always @(*) begin
        P1_P2_be3 = P1_P2_P3_BE_n; $display(";A 111");		//(= P1_P2_be3    P1_P2_P3_BE_n )) ;111
    end

    always @(*) begin
        P1_P2_addr3 = P1_P2_P3_Address; $display(";A 112");		//(= P1_P2_addr3    P1_P2_P3_Address )) ;112
    end

    always @(*) begin
        P1_P2_wr3 = P1_P2_P3_W_R_n; $display(";A 113");		//(= P1_P2_wr3    P1_P2_P3_W_R_n )) ;113
    end

    always @(*) begin
        P1_P2_dc3 = P1_P2_P3_D_C_n; $display(";A 114");		//(= P1_P2_dc3    P1_P2_P3_D_C_n )) ;114
    end

    always @(*) begin
        P1_P2_mio3 = P1_P2_P3_M_IO_n; $display(";A 115");		//(= P1_P2_mio3    P1_P2_P3_M_IO_n )) ;115
    end

    always @(*) begin
        P1_P2_ads3 = P1_P2_P3_ADS_n; $display(";A 116");		//(= P1_P2_ads3    P1_P2_P3_ADS_n )) ;116
    end

    always @(*) begin
        P1_P2_P3_Datai = P1_P2_di3; $display(";A 117");		//(= P1_P2_P3_Datai    P1_P2_di3 )) ;117
    end

    always @(*) begin
        P1_P2_do3 = P1_P2_P3_Datao; $display(";A 118");		//(= P1_P2_do3    P1_P2_P3_Datao )) ;118
    end

    always @(*) begin
        P1_P2_P3_CLOCK = P1_P2_clock; $display(";A 119");		//(= P1_P2_P3_CLOCK    P1_P2_clock )) ;119
    end

    always @(*) begin
        P1_P2_P3_NA_n = P1_P2_na; $display(";A 120");		//(= P1_P2_P3_NA_n    P1_P2_na )) ;120
    end

    always @(*) begin
        P1_P2_P3_BS16_n = P1_P2_bs16; $display(";A 121");		//(= P1_P2_P3_BS16_n    P1_P2_bs16 )) ;121
    end

    always @(*) begin
        P1_P2_P3_READY_n = P1_P2_rdy3; $display(";A 122");		//(= P1_P2_P3_READY_n    P1_P2_rdy3 )) ;122
    end

    always @(*) begin
        P1_P2_P3_HOLD = P1_P2_hold; $display(";A 123");		//(= P1_P2_P3_HOLD    P1_P2_hold )) ;123
    end

    always @(*) begin
        P1_P2_P3_RESET = P1_P2_reset;    end

    always @(*) begin
        P1_P3_clock = P1_clock; $display(";A 125");		//(= P1_P3_clock    P1_clock )) ;125
    end

    always @(*) begin
        P1_P3_reset = P1_reset;    end

    always @(*) begin
        P1_ad31 = P1_P3_addr; $display(";A 127");		//(= P1_ad31    P1_P3_addr )) ;127
    end

    always @(*) begin
        P1_P3_datai = P1_di3; $display(";A 128");		//(= P1_P3_datai    P1_di3 )) ;128
    end

    always @(*) begin
        P1_do3 = P1_P3_datao; $display(";A 129");		//(= P1_do3    P1_P3_datao )) ;129
    end

    always @(*) begin
        P1_rd3 = P1_P3_rd; $display(";A 130");		//(= P1_rd3    P1_P3_rd )) ;130
    end

    always @(*) begin
        P1_wr3 = P1_P3_wr; $display(";A 131");		//(= P1_wr3    P1_P3_wr )) ;131
    end

    always @(*) begin
        P1_P4_clock = P1_clock; $display(";A 132");		//(= P1_P4_clock    P1_clock )) ;132
    end

    always @(*) begin
        P1_P4_reset = P1_reset;    end

    always @(*) begin
        P1_ad41 = P1_P4_addr; $display(";A 134");		//(= P1_ad41    P1_P4_addr )) ;134
    end

    always @(*) begin
        P1_P4_datai = P1_di4; $display(";A 135");		//(= P1_P4_datai    P1_di4 )) ;135
    end

    always @(*) begin
        P1_do4 = P1_P4_datao; $display(";A 136");		//(= P1_do4    P1_P4_datao )) ;136
    end

    always @(*) begin
        P1_rd4 = P1_P4_rd; $display(";A 137");		//(= P1_rd4    P1_P4_rd )) ;137
    end

    always @(*) begin
        P1_wr4 = P1_P4_wr; $display(";A 138");		//(= P1_wr4    P1_P4_wr )) ;138
    end

    always @(*) begin
        P2_clock = clock; $display(";A 139");		//(= P2_clock    clock )) ;139
    end

    always @(*) begin
        P2_reset = reset;    end

    always @(*) begin
        P2_hold = hold; $display(";A 141");		//(= P2_hold    hold )) ;141
    end

    always @(*) begin
        P2_na = na; $display(";A 142");		//(= P2_na    na )) ;142
    end

    always @(*) begin
        P2_bs = bs; $display(";A 143");		//(= P2_bs    bs )) ;143
    end

    always @(*) begin
        P2_sel = sel2; $display(";A 144");		//(= P2_sel    sel2 )) ;144
    end

    always @(*) begin
        do2 = P2_dout; $display(";A 145");		//(= do2    P2_dout )) ;145
    end

    always @(*) begin
        P2_din = di2; $display(";A 146");		//(= P2_din    di2 )) ;146
    end

    always @(*) begin
        ax2 = P2_aux; $display(";A 147");		//(= ax2    P2_aux )) ;147
    end

    always @(*) begin
        P2_P1_clock = P2_clock; $display(";A 148");		//(= P2_P1_clock    P2_clock )) ;148
    end

    always @(*) begin
        P2_P1_reset = P2_reset;    end

    always @(*) begin
        P2_P1_datai = P2_di1; $display(";A 150");		//(= P2_P1_datai    P2_di1 )) ;150
    end

    always @(*) begin
        P2_do1 = P2_P1_datao; $display(";A 151");		//(= P2_do1    P2_P1_datao )) ;151
    end

    always @(*) begin
        P2_P1_hold = P2_hold; $display(";A 152");		//(= P2_P1_hold    P2_hold )) ;152
    end

    always @(*) begin
        P2_P1_na = P2_na; $display(";A 153");		//(= P2_P1_na    P2_na )) ;153
    end

    always @(*) begin
        P2_P1_bs16 = P2_bs; $display(";A 154");		//(= P2_P1_bs16    P2_bs )) ;154
    end

    always @(*) begin
        P2_ad11 = P2_P1_address1; $display(";A 155");		//(= P2_ad11    P2_P1_address1 )) ;155
    end

    always @(*) begin
        P2_ad12 = P2_P1_address2; $display(";A 156");		//(= P2_ad12    P2_P1_address2 )) ;156
    end

    always @(*) begin
        P2_wr1 = P2_P1_wr; $display(";A 157");		//(= P2_wr1    P2_P1_wr )) ;157
    end

    always @(*) begin
        P2_dc1 = P2_P1_dc; $display(";A 158");		//(= P2_dc1    P2_P1_dc )) ;158
    end

    always @(*) begin
        P2_mio1 = P2_P1_mio; $display(";A 159");		//(= P2_mio1    P2_P1_mio )) ;159
    end

    always @(*) begin
        P2_as11 = P2_P1_ast1; $display(";A 160");		//(= P2_as11    P2_P1_ast1 )) ;160
    end

    always @(*) begin
        P2_as12 = P2_P1_ast2; $display(";A 161");		//(= P2_as12    P2_P1_ast2 )) ;161
    end

    always @(*) begin
        P2_P1_ready1 = P2_r11; $display(";A 162");		//(= P2_P1_ready1    P2_r11 )) ;162
    end

    always @(*) begin
        P2_P1_ready2 = P2_r12; $display(";A 163");		//(= P2_P1_ready2    P2_r12 )) ;163
    end

    always @(*) begin
        P2_P1_be1 = P2_P1_P1_BE_n; $display(";A 164");		//(= P2_P1_be1    P2_P1_P1_BE_n )) ;164
    end

    always @(*) begin
        P2_P1_addr1 = P2_P1_P1_Address; $display(";A 165");		//(= P2_P1_addr1    P2_P1_P1_Address )) ;165
    end

    always @(*) begin
        P2_P1_wr1 = P2_P1_P1_W_R_n; $display(";A 166");		//(= P2_P1_wr1    P2_P1_P1_W_R_n )) ;166
    end

    always @(*) begin
        P2_P1_dc1 = P2_P1_P1_D_C_n; $display(";A 167");		//(= P2_P1_dc1    P2_P1_P1_D_C_n )) ;167
    end

    always @(*) begin
        P2_P1_mio1 = P2_P1_P1_M_IO_n; $display(";A 168");		//(= P2_P1_mio1    P2_P1_P1_M_IO_n )) ;168
    end

    always @(*) begin
        P2_P1_ads1 = P2_P1_P1_ADS_n; $display(";A 169");		//(= P2_P1_ads1    P2_P1_P1_ADS_n )) ;169
    end

    always @(*) begin
        P2_P1_P1_Datai = P2_P1_di1; $display(";A 170");		//(= P2_P1_P1_Datai    P2_P1_di1 )) ;170
    end

    always @(*) begin
        P2_P1_do1 = P2_P1_P1_Datao; $display(";A 171");		//(= P2_P1_do1    P2_P1_P1_Datao )) ;171
    end

    always @(*) begin
        P2_P1_P1_CLOCK = P2_P1_clock; $display(";A 172");		//(= P2_P1_P1_CLOCK    P2_P1_clock )) ;172
    end

    always @(*) begin
        P2_P1_P1_NA_n = P2_P1_na; $display(";A 173");		//(= P2_P1_P1_NA_n    P2_P1_na )) ;173
    end

    always @(*) begin
        P2_P1_P1_BS16_n = P2_P1_bs16; $display(";A 174");		//(= P2_P1_P1_BS16_n    P2_P1_bs16 )) ;174
    end

    always @(*) begin
        P2_P1_P1_READY_n = P2_P1_rdy1; $display(";A 175");		//(= P2_P1_P1_READY_n    P2_P1_rdy1 )) ;175
    end

    always @(*) begin
        P2_P1_P1_HOLD = P2_P1_hold; $display(";A 176");		//(= P2_P1_P1_HOLD    P2_P1_hold )) ;176
    end

    always @(*) begin
        P2_P1_P1_RESET = P2_P1_reset;    end

    always @(*) begin
        P2_P1_be2 = P2_P1_P2_BE_n; $display(";A 178");		//(= P2_P1_be2    P2_P1_P2_BE_n )) ;178
    end

    always @(*) begin
        P2_P1_addr2 = P2_P1_P2_Address; $display(";A 179");		//(= P2_P1_addr2    P2_P1_P2_Address )) ;179
    end

    always @(*) begin
        P2_P1_wr2 = P2_P1_P2_W_R_n; $display(";A 180");		//(= P2_P1_wr2    P2_P1_P2_W_R_n )) ;180
    end

    always @(*) begin
        P2_P1_dc2 = P2_P1_P2_D_C_n; $display(";A 181");		//(= P2_P1_dc2    P2_P1_P2_D_C_n )) ;181
    end

    always @(*) begin
        P2_P1_mio2 = P2_P1_P2_M_IO_n; $display(";A 182");		//(= P2_P1_mio2    P2_P1_P2_M_IO_n )) ;182
    end

    always @(*) begin
        P2_P1_ads2 = P2_P1_P2_ADS_n; $display(";A 183");		//(= P2_P1_ads2    P2_P1_P2_ADS_n )) ;183
    end

    always @(*) begin
        P2_P1_P2_Datai = P2_P1_di2; $display(";A 184");		//(= P2_P1_P2_Datai    P2_P1_di2 )) ;184
    end

    always @(*) begin
        P2_P1_do2 = P2_P1_P2_Datao; $display(";A 185");		//(= P2_P1_do2    P2_P1_P2_Datao )) ;185
    end

    always @(*) begin
        P2_P1_P2_CLOCK = P2_P1_clock; $display(";A 186");		//(= P2_P1_P2_CLOCK    P2_P1_clock )) ;186
    end

    always @(*) begin
        P2_P1_P2_NA_n = P2_P1_na; $display(";A 187");		//(= P2_P1_P2_NA_n    P2_P1_na )) ;187
    end

    always @(*) begin
        P2_P1_P2_BS16_n = P2_P1_bs16; $display(";A 188");		//(= P2_P1_P2_BS16_n    P2_P1_bs16 )) ;188
    end

    always @(*) begin
        P2_P1_P2_READY_n = P2_P1_rdy2; $display(";A 189");		//(= P2_P1_P2_READY_n    P2_P1_rdy2 )) ;189
    end

    always @(*) begin
        P2_P1_P2_HOLD = P2_P1_hold; $display(";A 190");		//(= P2_P1_P2_HOLD    P2_P1_hold )) ;190
    end

    always @(*) begin
        P2_P1_P2_RESET = P2_P1_reset;    end

    always @(*) begin
        P2_P1_be3 = P2_P1_P3_BE_n; $display(";A 192");		//(= P2_P1_be3    P2_P1_P3_BE_n )) ;192
    end

    always @(*) begin
        P2_P1_addr3 = P2_P1_P3_Address; $display(";A 193");		//(= P2_P1_addr3    P2_P1_P3_Address )) ;193
    end

    always @(*) begin
        P2_P1_wr3 = P2_P1_P3_W_R_n; $display(";A 194");		//(= P2_P1_wr3    P2_P1_P3_W_R_n )) ;194
    end

    always @(*) begin
        P2_P1_dc3 = P2_P1_P3_D_C_n; $display(";A 195");		//(= P2_P1_dc3    P2_P1_P3_D_C_n )) ;195
    end

    always @(*) begin
        P2_P1_mio3 = P2_P1_P3_M_IO_n; $display(";A 196");		//(= P2_P1_mio3    P2_P1_P3_M_IO_n )) ;196
    end

    always @(*) begin
        P2_P1_ads3 = P2_P1_P3_ADS_n; $display(";A 197");		//(= P2_P1_ads3    P2_P1_P3_ADS_n )) ;197
    end

    always @(*) begin
        P2_P1_P3_Datai = P2_P1_di3; $display(";A 198");		//(= P2_P1_P3_Datai    P2_P1_di3 )) ;198
    end

    always @(*) begin
        P2_P1_do3 = P2_P1_P3_Datao; $display(";A 199");		//(= P2_P1_do3    P2_P1_P3_Datao )) ;199
    end

    always @(*) begin
        P2_P1_P3_CLOCK = P2_P1_clock; $display(";A 200");		//(= P2_P1_P3_CLOCK    P2_P1_clock )) ;200
    end

    always @(*) begin
        P2_P1_P3_NA_n = P2_P1_na; $display(";A 201");		//(= P2_P1_P3_NA_n    P2_P1_na )) ;201
    end

    always @(*) begin
        P2_P1_P3_BS16_n = P2_P1_bs16; $display(";A 202");		//(= P2_P1_P3_BS16_n    P2_P1_bs16 )) ;202
    end

    always @(*) begin
        P2_P1_P3_READY_n = P2_P1_rdy3; $display(";A 203");		//(= P2_P1_P3_READY_n    P2_P1_rdy3 )) ;203
    end

    always @(*) begin
        P2_P1_P3_HOLD = P2_P1_hold; $display(";A 204");		//(= P2_P1_P3_HOLD    P2_P1_hold )) ;204
    end

    always @(*) begin
        P2_P1_P3_RESET = P2_P1_reset;    end

    always @(*) begin
        P2_P2_clock = P2_clock; $display(";A 206");		//(= P2_P2_clock    P2_clock )) ;206
    end

    always @(*) begin
        P2_P2_reset = P2_reset;    end

    always @(*) begin
        P2_P2_datai = P2_di2; $display(";A 208");		//(= P2_P2_datai    P2_di2 )) ;208
    end

    always @(*) begin
        P2_do2 = P2_P2_datao; $display(";A 209");		//(= P2_do2    P2_P2_datao )) ;209
    end

    always @(*) begin
        P2_P2_hold = P2_hold; $display(";A 210");		//(= P2_P2_hold    P2_hold )) ;210
    end

    always @(*) begin
        P2_P2_na = P2_na; $display(";A 211");		//(= P2_P2_na    P2_na )) ;211
    end

    always @(*) begin
        P2_P2_bs16 = P2_bs; $display(";A 212");		//(= P2_P2_bs16    P2_bs )) ;212
    end

    always @(*) begin
        P2_ad21 = P2_P2_address1; $display(";A 213");		//(= P2_ad21    P2_P2_address1 )) ;213
    end

    always @(*) begin
        P2_ad22 = P2_P2_address2; $display(";A 214");		//(= P2_ad22    P2_P2_address2 )) ;214
    end

    always @(*) begin
        P2_wr2 = P2_P2_wr; $display(";A 215");		//(= P2_wr2    P2_P2_wr )) ;215
    end

    always @(*) begin
        P2_dc2 = P2_P2_dc; $display(";A 216");		//(= P2_dc2    P2_P2_dc )) ;216
    end

    always @(*) begin
        P2_mio2 = P2_P2_mio; $display(";A 217");		//(= P2_mio2    P2_P2_mio )) ;217
    end

    always @(*) begin
        P2_as21 = P2_P2_ast1; $display(";A 218");		//(= P2_as21    P2_P2_ast1 )) ;218
    end

    always @(*) begin
        P2_as22 = P2_P2_ast2; $display(";A 219");		//(= P2_as22    P2_P2_ast2 )) ;219
    end

    always @(*) begin
        P2_P2_ready1 = P2_r21; $display(";A 220");		//(= P2_P2_ready1    P2_r21 )) ;220
    end

    always @(*) begin
        P2_P2_ready2 = P2_r22; $display(";A 221");		//(= P2_P2_ready2    P2_r22 )) ;221
    end

    always @(*) begin
        P2_P2_be1 = P2_P2_P1_BE_n; $display(";A 222");		//(= P2_P2_be1    P2_P2_P1_BE_n )) ;222
    end

    always @(*) begin
        P2_P2_addr1 = P2_P2_P1_Address; $display(";A 223");		//(= P2_P2_addr1    P2_P2_P1_Address )) ;223
    end

    always @(*) begin
        P2_P2_wr1 = P2_P2_P1_W_R_n; $display(";A 224");		//(= P2_P2_wr1    P2_P2_P1_W_R_n )) ;224
    end

    always @(*) begin
        P2_P2_dc1 = P2_P2_P1_D_C_n; $display(";A 225");		//(= P2_P2_dc1    P2_P2_P1_D_C_n )) ;225
    end

    always @(*) begin
        P2_P2_mio1 = P2_P2_P1_M_IO_n; $display(";A 226");		//(= P2_P2_mio1    P2_P2_P1_M_IO_n )) ;226
    end

    always @(*) begin
        P2_P2_ads1 = P2_P2_P1_ADS_n; $display(";A 227");		//(= P2_P2_ads1    P2_P2_P1_ADS_n )) ;227
    end

    always @(*) begin
        P2_P2_P1_Datai = P2_P2_di1; $display(";A 228");		//(= P2_P2_P1_Datai    P2_P2_di1 )) ;228
    end

    always @(*) begin
        P2_P2_do1 = P2_P2_P1_Datao; $display(";A 229");		//(= P2_P2_do1    P2_P2_P1_Datao )) ;229
    end

    always @(*) begin
        P2_P2_P1_CLOCK = P2_P2_clock; $display(";A 230");		//(= P2_P2_P1_CLOCK    P2_P2_clock )) ;230
    end

    always @(*) begin
        P2_P2_P1_NA_n = P2_P2_na; $display(";A 231");		//(= P2_P2_P1_NA_n    P2_P2_na )) ;231
    end

    always @(*) begin
        P2_P2_P1_BS16_n = P2_P2_bs16; $display(";A 232");		//(= P2_P2_P1_BS16_n    P2_P2_bs16 )) ;232
    end

    always @(*) begin
        P2_P2_P1_READY_n = P2_P2_rdy1; $display(";A 233");		//(= P2_P2_P1_READY_n    P2_P2_rdy1 )) ;233
    end

    always @(*) begin
        P2_P2_P1_HOLD = P2_P2_hold; $display(";A 234");		//(= P2_P2_P1_HOLD    P2_P2_hold )) ;234
    end

    always @(*) begin
        P2_P2_P1_RESET = P2_P2_reset;    end

    always @(*) begin
        P2_P2_be2 = P2_P2_P2_BE_n; $display(";A 236");		//(= P2_P2_be2    P2_P2_P2_BE_n )) ;236
    end

    always @(*) begin
        P2_P2_addr2 = P2_P2_P2_Address; $display(";A 237");		//(= P2_P2_addr2    P2_P2_P2_Address )) ;237
    end

    always @(*) begin
        P2_P2_wr2 = P2_P2_P2_W_R_n; $display(";A 238");		//(= P2_P2_wr2    P2_P2_P2_W_R_n )) ;238
    end

    always @(*) begin
        P2_P2_dc2 = P2_P2_P2_D_C_n; $display(";A 239");		//(= P2_P2_dc2    P2_P2_P2_D_C_n )) ;239
    end

    always @(*) begin
        P2_P2_mio2 = P2_P2_P2_M_IO_n; $display(";A 240");		//(= P2_P2_mio2    P2_P2_P2_M_IO_n )) ;240
    end

    always @(*) begin
        P2_P2_ads2 = P2_P2_P2_ADS_n; $display(";A 241");		//(= P2_P2_ads2    P2_P2_P2_ADS_n )) ;241
    end

    always @(*) begin
        P2_P2_P2_Datai = P2_P2_di2; $display(";A 242");		//(= P2_P2_P2_Datai    P2_P2_di2 )) ;242
    end

    always @(*) begin
        P2_P2_do2 = P2_P2_P2_Datao; $display(";A 243");		//(= P2_P2_do2    P2_P2_P2_Datao )) ;243
    end

    always @(*) begin
        P2_P2_P2_CLOCK = P2_P2_clock; $display(";A 244");		//(= P2_P2_P2_CLOCK    P2_P2_clock )) ;244
    end

    always @(*) begin
        P2_P2_P2_NA_n = P2_P2_na; $display(";A 245");		//(= P2_P2_P2_NA_n    P2_P2_na )) ;245
    end

    always @(*) begin
        P2_P2_P2_BS16_n = P2_P2_bs16; $display(";A 246");		//(= P2_P2_P2_BS16_n    P2_P2_bs16 )) ;246
    end

    always @(*) begin
        P2_P2_P2_READY_n = P2_P2_rdy2; $display(";A 247");		//(= P2_P2_P2_READY_n    P2_P2_rdy2 )) ;247
    end

    always @(*) begin
        P2_P2_P2_HOLD = P2_P2_hold; $display(";A 248");		//(= P2_P2_P2_HOLD    P2_P2_hold )) ;248
    end

    always @(*) begin
        P2_P2_P2_RESET = P2_P2_reset;    end

    always @(*) begin
        P2_P2_be3 = P2_P2_P3_BE_n; $display(";A 250");		//(= P2_P2_be3    P2_P2_P3_BE_n )) ;250
    end

    always @(*) begin
        P2_P2_addr3 = P2_P2_P3_Address; $display(";A 251");		//(= P2_P2_addr3    P2_P2_P3_Address )) ;251
    end

    always @(*) begin
        P2_P2_wr3 = P2_P2_P3_W_R_n; $display(";A 252");		//(= P2_P2_wr3    P2_P2_P3_W_R_n )) ;252
    end

    always @(*) begin
        P2_P2_dc3 = P2_P2_P3_D_C_n; $display(";A 253");		//(= P2_P2_dc3    P2_P2_P3_D_C_n )) ;253
    end

    always @(*) begin
        P2_P2_mio3 = P2_P2_P3_M_IO_n; $display(";A 254");		//(= P2_P2_mio3    P2_P2_P3_M_IO_n )) ;254
    end

    always @(*) begin
        P2_P2_ads3 = P2_P2_P3_ADS_n; $display(";A 255");		//(= P2_P2_ads3    P2_P2_P3_ADS_n )) ;255
    end

    always @(*) begin
        P2_P2_P3_Datai = P2_P2_di3; $display(";A 256");		//(= P2_P2_P3_Datai    P2_P2_di3 )) ;256
    end

    always @(*) begin
        P2_P2_do3 = P2_P2_P3_Datao; $display(";A 257");		//(= P2_P2_do3    P2_P2_P3_Datao )) ;257
    end

    always @(*) begin
        P2_P2_P3_CLOCK = P2_P2_clock; $display(";A 258");		//(= P2_P2_P3_CLOCK    P2_P2_clock )) ;258
    end

    always @(*) begin
        P2_P2_P3_NA_n = P2_P2_na; $display(";A 259");		//(= P2_P2_P3_NA_n    P2_P2_na )) ;259
    end

    always @(*) begin
        P2_P2_P3_BS16_n = P2_P2_bs16; $display(";A 260");		//(= P2_P2_P3_BS16_n    P2_P2_bs16 )) ;260
    end

    always @(*) begin
        P2_P2_P3_READY_n = P2_P2_rdy3; $display(";A 261");		//(= P2_P2_P3_READY_n    P2_P2_rdy3 )) ;261
    end

    always @(*) begin
        P2_P2_P3_HOLD = P2_P2_hold; $display(";A 262");		//(= P2_P2_P3_HOLD    P2_P2_hold )) ;262
    end

    always @(*) begin
        P2_P2_P3_RESET = P2_P2_reset;    end

    always @(*) begin
        P2_P3_clock = P2_clock; $display(";A 264");		//(= P2_P3_clock    P2_clock )) ;264
    end

    always @(*) begin
        P2_P3_reset = P2_reset;    end

    always @(*) begin
        P2_ad31 = P2_P3_addr; $display(";A 266");		//(= P2_ad31    P2_P3_addr )) ;266
    end

    always @(*) begin
        P2_P3_datai = P2_di3; $display(";A 267");		//(= P2_P3_datai    P2_di3 )) ;267
    end

    always @(*) begin
        P2_do3 = P2_P3_datao; $display(";A 268");		//(= P2_do3    P2_P3_datao )) ;268
    end

    always @(*) begin
        P2_rd3 = P2_P3_rd; $display(";A 269");		//(= P2_rd3    P2_P3_rd )) ;269
    end

    always @(*) begin
        P2_wr3 = P2_P3_wr; $display(";A 270");		//(= P2_wr3    P2_P3_wr )) ;270
    end

    always @(*) begin
        P2_P4_clock = P2_clock; $display(";A 271");		//(= P2_P4_clock    P2_clock )) ;271
    end

    always @(*) begin
        P2_P4_reset = P2_reset;    end

    always @(*) begin
        P2_ad41 = P2_P4_addr; $display(";A 273");		//(= P2_ad41    P2_P4_addr )) ;273
    end

    always @(*) begin
        P2_P4_datai = P2_di4; $display(";A 274");		//(= P2_P4_datai    P2_di4 )) ;274
    end

    always @(*) begin
        P2_do4 = P2_P4_datao; $display(";A 275");		//(= P2_do4    P2_P4_datao )) ;275
    end

    always @(*) begin
        P2_rd4 = P2_P4_rd; $display(";A 276");		//(= P2_rd4    P2_P4_rd )) ;276
    end

    always @(*) begin
        P2_wr4 = P2_P4_wr; $display(";A 277");		//(= P2_wr4    P2_P4_wr )) ;277
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:144
    always @(posedge P1_P1_reset or posedge P1_P1_clock) begin
        if ((P1_P1_reset == 1'b1)) begin
            P1_P1_buf1 <= #1 32'sb00000000000000000000000000000000; $display(";A 280");		//(= P1_P1_buf1    0b00000000000000000000000000000000)) ;280
            P1_P1_ready11 <= #1 1'b0; $display(";A 281");		//(= P1_P1_ready11    0b0)) ;281
            P1_P1_ready12 <= #1 1'b0; $display(";A 282");		//(= P1_P1_ready12    0b0)) ;282
        end
        else begin
            if (((((((P1_P1_addr1 > 30'b100000000000000000000000000000) & (P1_P1_ads1 == 1'b0)) & (P1_P1_mio1 == 1'b1)) & (P1_P1_dc1 == 1'b0)) & (P1_P1_wr1 == 1'b1)) & (P1_P1_be1 == 4'b0000))) begin
                $display(";A 283");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P1_addr1  0b100000000000000000000000000000)) (bv-comp P1_P1_ads1  0b0)) (bv-comp P1_P1_mio1  0b1)) (bv-comp P1_P1_dc1  0b0)) (bv-comp P1_P1_wr1  0b1)) (bv-comp P1_P1_be1  0b0000))   0b1)) ;283
                P1_P1_buf1 <= #1 P1_P1_do1; $display(";A 285");		//(= P1_P1_buf1    P1_P1_do1 )) ;285
                P1_P1_ready11 <= #1 1'b0; $display(";A 286");		//(= P1_P1_ready11    0b0)) ;286
                P1_P1_ready12 <= #1 1'b1; $display(";A 287");		//(= P1_P1_ready12    0b1)) ;287
            end
            else begin
                $display(";A 284");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P1_addr1  0b100000000000000000000000000000)) (bv-comp P1_P1_ads1  0b0)) (bv-comp P1_P1_mio1  0b1)) (bv-comp P1_P1_dc1  0b0)) (bv-comp P1_P1_wr1  0b1)) (bv-comp P1_P1_be1  0b0000))   0b0)) ;284
                if (((((((P1_P1_addr2 > 30'b100000000000000000000000000000) & (P1_P1_ads2 == 1'b0)) & (P1_P1_mio2 == 1'b1)) & (P1_P1_dc2 == 1'b0)) & (P1_P1_wr2 == 1'b1)) & (P1_P1_be2 == 4'b0000))) begin
                    $display(";A 288");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P1_addr2  0b100000000000000000000000000000)) (bv-comp P1_P1_ads2  0b0)) (bv-comp P1_P1_mio2  0b1)) (bv-comp P1_P1_dc2  0b0)) (bv-comp P1_P1_wr2  0b1)) (bv-comp P1_P1_be2  0b0000))   0b1)) ;288
                    P1_P1_buf1 <= #1 P1_P1_do2; $display(";A 290");		//(= P1_P1_buf1    P1_P1_do2 )) ;290
                    P1_P1_ready11 <= #1 1'b1; $display(";A 291");		//(= P1_P1_ready11    0b1)) ;291
                    P1_P1_ready12 <= #1 1'b0; $display(";A 292");		//(= P1_P1_ready12    0b0)) ;292
                end
                else begin
                    $display(";A 289");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P1_addr2  0b100000000000000000000000000000)) (bv-comp P1_P1_ads2  0b0)) (bv-comp P1_P1_mio2  0b1)) (bv-comp P1_P1_dc2  0b0)) (bv-comp P1_P1_wr2  0b1)) (bv-comp P1_P1_be2  0b0000))   0b0)) ;289
                    P1_P1_ready11 <= #1 1'b1; $display(";A 293");		//(= P1_P1_ready11    0b1)) ;293
                    P1_P1_ready12 <= #1 1'b1; $display(";A 294");		//(= P1_P1_ready12    0b1)) ;294
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:173
    always @(posedge P1_P1_reset or posedge P1_P1_clock) begin
        if ((P1_P1_reset == 1'b1)) begin
            P1_P1_buf2 <= #1 32'sb00000000000000000000000000000000; $display(";A 297");		//(= P1_P1_buf2    0b00000000000000000000000000000000)) ;297
            P1_P1_ready21 <= #1 1'b0; $display(";A 298");		//(= P1_P1_ready21    0b0)) ;298
            P1_P1_ready22 <= #1 1'b0; $display(";A 299");		//(= P1_P1_ready22    0b0)) ;299
        end
        else begin
            if (((((((P1_P1_addr2 < 30'b100000000000000000000000000000) & (P1_P1_ads2 == 1'b0)) & (P1_P1_mio2 == 1'b1)) & (P1_P1_dc2 == 1'b0)) & (P1_P1_wr2 == 1'b1)) & (P1_P1_be2 == 4'b0000))) begin
                $display(";A 300");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P1_P1_addr2  0b100000000000000000000000000000)) (bv-comp P1_P1_ads2  0b0)) (bv-comp P1_P1_mio2  0b1)) (bv-comp P1_P1_dc2  0b0)) (bv-comp P1_P1_wr2  0b1)) (bv-comp P1_P1_be2  0b0000))   0b1)) ;300
                P1_P1_buf2 <= #1 P1_P1_do2; $display(";A 302");		//(= P1_P1_buf2    P1_P1_do2 )) ;302
                P1_P1_ready21 <= #1 1'b0; $display(";A 303");		//(= P1_P1_ready21    0b0)) ;303
                P1_P1_ready22 <= #1 1'b1; $display(";A 304");		//(= P1_P1_ready22    0b1)) ;304
            end
            else begin
                $display(";A 301");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P1_P1_addr2  0b100000000000000000000000000000)) (bv-comp P1_P1_ads2  0b0)) (bv-comp P1_P1_mio2  0b1)) (bv-comp P1_P1_dc2  0b0)) (bv-comp P1_P1_wr2  0b1)) (bv-comp P1_P1_be2  0b0000))   0b0)) ;301
                if ((((((P1_P1_ads3 == 1'b0) & (P1_P1_mio3 == 1'b1)) & (P1_P1_dc3 == 1'b0)) & (P1_P1_wr3 == 1'b0)) & (P1_P1_be3 == 4'b0000))) begin
                    $display(";A 305");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P1_P1_ads3  0b0) (bv-comp P1_P1_mio3  0b1)) (bv-comp P1_P1_dc3  0b0)) (bv-comp P1_P1_wr3  0b0)) (bv-comp P1_P1_be3  0b0000))   0b1)) ;305
                    P1_P1_ready21 <= #1 1'b1; $display(";A 307");		//(= P1_P1_ready21    0b1)) ;307
                    P1_P1_ready22 <= #1 1'b0; $display(";A 308");		//(= P1_P1_ready22    0b0)) ;308
                end
                else begin
                    $display(";A 306");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P1_P1_ads3  0b0) (bv-comp P1_P1_mio3  0b1)) (bv-comp P1_P1_dc3  0b0)) (bv-comp P1_P1_wr3  0b0)) (bv-comp P1_P1_be3  0b0000))   0b0)) ;306
                    P1_P1_ready21 <= #1 1'b1; $display(";A 309");		//(= P1_P1_ready21    0b1)) ;309
                    P1_P1_ready22 <= #1 1'b1; $display(";A 310");		//(= P1_P1_ready22    0b1)) ;310
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:201
    always @(P1_P1_datai or P1_P1_buf1 or P1_P1_addr1) begin
        if ((P1_P1_addr1 > 30'b100000000000000000000000000000)) begin
            $display(";A 311");		//(= (bool-to-bv (bv-gt P1_P1_addr1  0b100000000000000000000000000000))   0b1)) ;311
            P1_P1_di1 <= #1 P1_P1_buf1; $display(";A 313");		//(= P1_P1_di1    P1_P1_buf1 )) ;313
        end
        else begin
            $display(";A 312");		//(= (bool-to-bv (bv-gt P1_P1_addr1  0b100000000000000000000000000000))   0b0)) ;312
            P1_P1_di1 <= #1 P1_P1_datai; $display(";A 314");		//(= P1_P1_di1    P1_P1_datai )) ;314
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:207
    always @(P1_P1_buf2 or P1_P1_buf1 or P1_P1_addr2) begin
        if ((P1_P1_addr2 > 30'b100000000000000000000000000000)) begin
            $display(";A 315");		//(= (bool-to-bv (bv-gt P1_P1_addr2  0b100000000000000000000000000000))   0b1)) ;315
            P1_P1_di2 <= #1 P1_P1_buf1; $display(";A 317");		//(= P1_P1_di2    P1_P1_buf1 )) ;317
        end
        else begin
            $display(";A 316");		//(= (bool-to-bv (bv-gt P1_P1_addr2  0b100000000000000000000000000000))   0b0)) ;316
            P1_P1_di2 <= #1 P1_P1_buf2; $display(";A 318");		//(= P1_P1_di2    P1_P1_buf2 )) ;318
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:213
    always @(P1_P1_do3 or P1_P1_do2 or P1_P1_do1 or P1_P1_addr3 or P1_P1_addr2) begin
        if ((((P1_P1_do1 < 32'b00000000000000000000000000000000) & (P1_P1_do2 < 32'b00000000000000000000000000000000)) & (P1_P1_do3 < 32'b00000000000000000000000000000000))) begin
            $display(";A 319");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P1_P1_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P1_P1_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P1_P1_do3  0b00000000000000000000000000000000)))   0b1)) ;319
            P1_P1_address2 <= #1 P1_P1_addr3; $display(";A 321");		//(= P1_P1_address2    P1_P1_addr3 )) ;321
        end
        else begin
            $display(";A 320");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P1_P1_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P1_P1_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P1_P1_do3  0b00000000000000000000000000000000)))   0b0)) ;320
            P1_P1_address2 <= #1 P1_P1_addr2; $display(";A 322");		//(= P1_P1_address2    P1_P1_addr2 )) ;322
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:219
    always @(P1_P1_ready22 or P1_P1_ready21 or P1_P1_ready12 or P1_P1_ready11 or P1_P1_ready2 or P1_P1_ready1 or P1_P1_ads3 or P1_P1_ads1 or P1_P1_mio3 or P1_P1_dc3 or P1_P1_wr3 or P1_P1_addr1 or P1_P1_do3 or P1_P1_buf2) begin
        P1_P1_di3 <= #1 P1_P1_buf2; $display(";A 323");		//(= P1_P1_di3    P1_P1_buf2 )) ;323
        P1_P1_datao <= #1 P1_P1_do3; $display(";A 324");		//(= P1_P1_datao    P1_P1_do3 )) ;324
        P1_P1_address1 <= #1 P1_P1_addr1; $display(";A 325");		//(= P1_P1_address1    P1_P1_addr1 )) ;325
        P1_P1_wr <= #1 P1_P1_wr3; $display(";A 326");		//(= P1_P1_wr    P1_P1_wr3 )) ;326
        P1_P1_dc <= #1 P1_P1_dc3; $display(";A 327");		//(= P1_P1_dc    P1_P1_dc3 )) ;327
        P1_P1_mio <= #1 P1_P1_mio3; $display(";A 328");		//(= P1_P1_mio    P1_P1_mio3 )) ;328
        P1_P1_ast1 <= #1 P1_P1_ads1; $display(";A 329");		//(= P1_P1_ast1    P1_P1_ads1 )) ;329
        P1_P1_ast2 <= #1 P1_P1_ads3; $display(";A 330");		//(= P1_P1_ast2    P1_P1_ads3 )) ;330
        P1_P1_rdy1 <= #1 (P1_P1_ready11 & P1_P1_ready1); $display(";A 331");		//(= P1_P1_rdy1    (bv-and P1_P1_ready11  P1_P1_ready1 ))) ;331
        P1_P1_rdy2 <= #1 (P1_P1_ready12 & P1_P1_ready21); $display(";A 332");		//(= P1_P1_rdy2    (bv-and P1_P1_ready12  P1_P1_ready21 ))) ;332
        P1_P1_rdy3 <= #1 (P1_P1_ready22 & P1_P1_ready2); $display(";A 333");		//(= P1_P1_rdy3    (bv-and P1_P1_ready22  P1_P1_ready2 ))) ;333
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:344
    always @(posedge P1_P1_P1_RESET or posedge P1_P1_P1_CLOCK) begin
        if ((P1_P1_P1_RESET == 1'b1)) begin
            $display(";A 334");		//(= (bv-comp P1_P1_P1_RESET  0b1)   0b1)) ;334
            P1_P1_P1_BE_n <= #1 4'b0000; $display(";A 336");		//(= P1_P1_P1_BE_n    0b0000)) ;336
            P1_P1_P1_Address <= #1 30'sb000000000000000000000000000000; $display(";A 337");		//(= P1_P1_P1_Address    0b000000000000000000000000000000)) ;337
            P1_P1_P1_W_R_n <= #1 1'b0; $display(";A 338");		//(= P1_P1_P1_W_R_n    0b0)) ;338
            P1_P1_P1_D_C_n <= #1 1'b0; $display(";A 339");		//(= P1_P1_P1_D_C_n    0b0)) ;339
            P1_P1_P1_M_IO_n <= #1 1'b0; $display(";A 340");		//(= P1_P1_P1_M_IO_n    0b0)) ;340
            P1_P1_P1_ADS_n <= #1 1'b0; $display(";A 341");		//(= P1_P1_P1_ADS_n    0b0)) ;341
            P1_P1_P1_State <= #1 3'sb000; $display(";A 342");		//(= P1_P1_P1_State    0b000)) ;342
            P1_P1_P1_StateNA <= #1 1'b0; $display(";A 343");		//(= P1_P1_P1_StateNA    0b0)) ;343
            P1_P1_P1_StateBS16 <= #1 1'b0; $display(";A 344");		//(= P1_P1_P1_StateBS16    0b0)) ;344
            P1_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 345");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000000)) ;345
        end
        else begin
            $display(";A 335");		//(= (bv-comp P1_P1_P1_RESET  0b1)   0b0)) ;335
            case (P1_P1_P1_State)
                3'b000 :
                    begin
                        $display(";A 346");		//(= P1_P1_P1_State    0b000)) ;346
                        P1_P1_P1_D_C_n <= #1 1'b1; $display(";A 347");		//(= P1_P1_P1_D_C_n    0b1)) ;347
                        P1_P1_P1_ADS_n <= #1 1'b1; $display(";A 348");		//(= P1_P1_P1_ADS_n    0b1)) ;348
                        P1_P1_P1_State <= #1 3'sb001; $display(";A 349");		//(= P1_P1_P1_State    0b001)) ;349
                        P1_P1_P1_StateNA <= #1 1'b1; $display(";A 350");		//(= P1_P1_P1_StateNA    0b1)) ;350
                        P1_P1_P1_StateBS16 <= #1 1'b1; $display(";A 351");		//(= P1_P1_P1_StateBS16    0b1)) ;351
                        P1_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 352");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;352
                        P1_P1_P1_State <= #1 3'sb001; $display(";A 353");		//(= P1_P1_P1_State    0b001)) ;353
                    end
                3'b001 :
                    begin
                        $display(";A 354");		//(= P1_P1_P1_State    0b001)) ;354
                        if ((P1_P1_P1_RequestPending == 1'b1)) begin
                            $display(";A 355");		//(= (bv-comp P1_P1_P1_RequestPending  0b1)   0b1)) ;355
                            P1_P1_P1_State <= #1 3'sb010; $display(";A 357");		//(= P1_P1_P1_State    0b010)) ;357
                        end
                        else begin
                            $display(";A 356");		//(= (bv-comp P1_P1_P1_RequestPending  0b1)   0b0)) ;356
                            if ((P1_P1_P1_HOLD == 1'b1)) begin
                                $display(";A 358");		//(= (bv-comp P1_P1_P1_HOLD  0b1)   0b1)) ;358
                                P1_P1_P1_State <= #1 3'sb101; $display(";A 360");		//(= P1_P1_P1_State    0b101)) ;360
                            end
                            else begin
                                $display(";A 359");		//(= (bv-comp P1_P1_P1_HOLD  0b1)   0b0)) ;359
                                P1_P1_P1_State <= #1 3'sb001; $display(";A 361");		//(= P1_P1_P1_State    0b001)) ;361
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 362");		//(= P1_P1_P1_State    0b010)) ;362
                        P1_P1_P1_Address <= #1 ((P1_P1_P1_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 363");		//(= P1_P1_P1_Address    (bv-smod (bv-sdiv P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;363
                        P1_P1_P1_BE_n <= #1 P1_P1_P1_ByteEnable; $display(";A 364");		//(= P1_P1_P1_BE_n    P1_P1_P1_ByteEnable )) ;364
                        P1_P1_P1_M_IO_n <= #1 P1_P1_P1_MemoryFetch; $display(";A 365");		//(= P1_P1_P1_M_IO_n    P1_P1_P1_MemoryFetch )) ;365
                        if ((P1_P1_P1_ReadRequest == 1'b1)) begin
                            $display(";A 366");		//(= (bv-comp P1_P1_P1_ReadRequest  0b1)   0b1)) ;366
                            P1_P1_P1_W_R_n <= #1 1'b0; $display(";A 368");		//(= P1_P1_P1_W_R_n    0b0)) ;368
                        end
                        else begin
                            $display(";A 367");		//(= (bv-comp P1_P1_P1_ReadRequest  0b1)   0b0)) ;367
                            P1_P1_P1_W_R_n <= #1 1'b1; $display(";A 369");		//(= P1_P1_P1_W_R_n    0b1)) ;369
                        end
                        if ((P1_P1_P1_CodeFetch == 1'b1)) begin
                            $display(";A 370");		//(= (bv-comp P1_P1_P1_CodeFetch  0b1)   0b1)) ;370
                            P1_P1_P1_D_C_n <= #1 1'b0; $display(";A 372");		//(= P1_P1_P1_D_C_n    0b0)) ;372
                        end
                        else begin
                            $display(";A 371");		//(= (bv-comp P1_P1_P1_CodeFetch  0b1)   0b0)) ;371
                            P1_P1_P1_D_C_n <= #1 1'b1; $display(";A 373");		//(= P1_P1_P1_D_C_n    0b1)) ;373
                        end
                        P1_P1_P1_ADS_n <= #1 1'b0; $display(";A 374");		//(= P1_P1_P1_ADS_n    0b0)) ;374
                        P1_P1_P1_State <= #1 3'sb011; $display(";A 375");		//(= P1_P1_P1_State    0b011)) ;375
                    end
                3'b011 :
                    begin
                        $display(";A 376");		//(= P1_P1_P1_State    0b011)) ;376
                        if ((((P1_P1_P1_READY_n == 1'b0) & (P1_P1_P1_HOLD == 1'b0)) & (P1_P1_P1_RequestPending == 1'b1))) begin
                            $display(";A 377");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b1))   0b1)) ;377
                            P1_P1_P1_State <= #1 3'sb010; $display(";A 379");		//(= P1_P1_P1_State    0b010)) ;379
                        end
                        else begin
                            $display(";A 378");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b1))   0b0)) ;378
                            if (((P1_P1_P1_READY_n == 1'b1) & (P1_P1_P1_NA_n == 1'b1))) begin
                                $display(";A 380");		//(= (bv-and (bv-comp P1_P1_P1_READY_n  0b1) (bv-comp P1_P1_P1_NA_n  0b1))   0b1)) ;380
                            end
                            else begin
                                $display(";A 381");		//(= (bv-and (bv-comp P1_P1_P1_READY_n  0b1) (bv-comp P1_P1_P1_NA_n  0b1))   0b0)) ;381
                                if ((((P1_P1_P1_RequestPending == 1'b1) | (P1_P1_P1_HOLD == 1'b1)) & ((P1_P1_P1_READY_n == 1'b1) & (P1_P1_P1_NA_n == 1'b0)))) begin
                                    $display(";A 382");		//(= (bv-and (bv-or (bv-comp P1_P1_P1_RequestPending  0b1) (bv-comp P1_P1_P1_HOLD  0b1)) (bv-and (bv-comp P1_P1_P1_READY_n  0b1) (bv-comp P1_P1_P1_NA_n  0b0)))   0b1)) ;382
                                    P1_P1_P1_State <= #1 3'sb111; $display(";A 384");		//(= P1_P1_P1_State    0b111)) ;384
                                end
                                else begin
                                    $display(";A 383");		//(= (bv-and (bv-or (bv-comp P1_P1_P1_RequestPending  0b1) (bv-comp P1_P1_P1_HOLD  0b1)) (bv-and (bv-comp P1_P1_P1_READY_n  0b1) (bv-comp P1_P1_P1_NA_n  0b0)))   0b0)) ;383
                                    if (((((P1_P1_P1_RequestPending == 1'b1) & (P1_P1_P1_HOLD == 1'b0)) & (P1_P1_P1_READY_n == 1'b1)) & (P1_P1_P1_NA_n == 1'b0))) begin
                                        $display(";A 385");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P1_P1_RequestPending  0b1) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_READY_n  0b1)) (bv-comp P1_P1_P1_NA_n  0b0))   0b1)) ;385
                                        P1_P1_P1_State <= #1 3'sb110; $display(";A 387");		//(= P1_P1_P1_State    0b110)) ;387
                                    end
                                    else begin
                                        $display(";A 386");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P1_P1_RequestPending  0b1) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_READY_n  0b1)) (bv-comp P1_P1_P1_NA_n  0b0))   0b0)) ;386
                                        if ((((P1_P1_P1_RequestPending == 1'b0) & (P1_P1_P1_HOLD == 1'b0)) & (P1_P1_P1_READY_n == 1'b0))) begin
                                            $display(";A 388");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_RequestPending  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_READY_n  0b0))   0b1)) ;388
                                            P1_P1_P1_State <= #1 3'sb001; $display(";A 390");		//(= P1_P1_P1_State    0b001)) ;390
                                        end
                                        else begin
                                            $display(";A 389");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_RequestPending  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_READY_n  0b0))   0b0)) ;389
                                            if (((P1_P1_P1_HOLD == 1'b1) & (P1_P1_P1_READY_n == 1'b1))) begin
                                                $display(";A 391");		//(= (bv-and (bv-comp P1_P1_P1_HOLD  0b1) (bv-comp P1_P1_P1_READY_n  0b1))   0b1)) ;391
                                                P1_P1_P1_State <= #1 3'sb101; $display(";A 393");		//(= P1_P1_P1_State    0b101)) ;393
                                            end
                                            else begin
                                                $display(";A 392");		//(= (bv-and (bv-comp P1_P1_P1_HOLD  0b1) (bv-comp P1_P1_P1_READY_n  0b1))   0b0)) ;392
                                                P1_P1_P1_State <= #1 3'sb011; $display(";A 394");		//(= P1_P1_P1_State    0b011)) ;394
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P1_P1_P1_StateBS16 <= #1 P1_P1_P1_BS16_n; $display(";A 395");		//(= P1_P1_P1_StateBS16    P1_P1_P1_BS16_n )) ;395
                        if ((P1_P1_P1_BS16_n == 1'b0)) begin
                            $display(";A 396");		//(= (bv-comp P1_P1_P1_BS16_n  0b0)   0b1)) ;396
                            P1_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 398");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000001)) ;398
                        end
                        else begin
                            $display(";A 397");		//(= (bv-comp P1_P1_P1_BS16_n  0b0)   0b0)) ;397
                            P1_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 399");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;399
                        end
                        P1_P1_P1_StateNA <= #1 P1_P1_P1_NA_n; $display(";A 400");		//(= P1_P1_P1_StateNA    P1_P1_P1_NA_n )) ;400
                        P1_P1_P1_ADS_n <= #1 1'b1; $display(";A 401");		//(= P1_P1_P1_ADS_n    0b1)) ;401
                    end
                3'b100 :
                    begin
                        $display(";A 402");		//(= P1_P1_P1_State    0b100)) ;402
                        if ((((P1_P1_P1_NA_n == 1'b0) & (P1_P1_P1_HOLD == 1'b0)) & (P1_P1_P1_RequestPending == 1'b1))) begin
                            $display(";A 403");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_NA_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b1))   0b1)) ;403
                            P1_P1_P1_State <= #1 3'sb110; $display(";A 405");		//(= P1_P1_P1_State    0b110)) ;405
                        end
                        else begin
                            $display(";A 404");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_NA_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b1))   0b0)) ;404
                            if (((P1_P1_P1_NA_n == 1'b0) & ((P1_P1_P1_HOLD == 1'b1) | (P1_P1_P1_RequestPending == 1'b0)))) begin
                                $display(";A 406");		//(= (bv-and (bv-comp P1_P1_P1_NA_n  0b0) (bv-or (bv-comp P1_P1_P1_HOLD  0b1) (bv-comp P1_P1_P1_RequestPending  0b0)))   0b1)) ;406
                                P1_P1_P1_State <= #1 3'sb111; $display(";A 408");		//(= P1_P1_P1_State    0b111)) ;408
                            end
                            else begin
                                $display(";A 407");		//(= (bv-and (bv-comp P1_P1_P1_NA_n  0b0) (bv-or (bv-comp P1_P1_P1_HOLD  0b1) (bv-comp P1_P1_P1_RequestPending  0b0)))   0b0)) ;407
                                if ((P1_P1_P1_NA_n == 1'b1)) begin
                                    $display(";A 409");		//(= (bv-comp P1_P1_P1_NA_n  0b1)   0b1)) ;409
                                    P1_P1_P1_State <= #1 3'sb011; $display(";A 411");		//(= P1_P1_P1_State    0b011)) ;411
                                end
                                else begin
                                    $display(";A 410");		//(= (bv-comp P1_P1_P1_NA_n  0b1)   0b0)) ;410
                                    P1_P1_P1_State <= #1 3'sb100; $display(";A 412");		//(= P1_P1_P1_State    0b100)) ;412
                                end
                            end
                        end
                        P1_P1_P1_StateBS16 <= #1 P1_P1_P1_BS16_n; $display(";A 413");		//(= P1_P1_P1_StateBS16    P1_P1_P1_BS16_n )) ;413
                        if ((P1_P1_P1_BS16_n == 1'b0)) begin
                            $display(";A 414");		//(= (bv-comp P1_P1_P1_BS16_n  0b0)   0b1)) ;414
                            P1_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 416");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000001)) ;416
                        end
                        else begin
                            $display(";A 415");		//(= (bv-comp P1_P1_P1_BS16_n  0b0)   0b0)) ;415
                            P1_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 417");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;417
                        end
                        P1_P1_P1_StateNA <= #1 P1_P1_P1_NA_n; $display(";A 418");		//(= P1_P1_P1_StateNA    P1_P1_P1_NA_n )) ;418
                        P1_P1_P1_ADS_n <= #1 1'b1; $display(";A 419");		//(= P1_P1_P1_ADS_n    0b1)) ;419
                    end
                3'b101 :
                    begin
                        $display(";A 420");		//(= P1_P1_P1_State    0b101)) ;420
                        if (((P1_P1_P1_HOLD == 1'b0) & (P1_P1_P1_RequestPending == 1'b1))) begin
                            $display(";A 421");		//(= (bv-and (bv-comp P1_P1_P1_HOLD  0b0) (bv-comp P1_P1_P1_RequestPending  0b1))   0b1)) ;421
                            P1_P1_P1_State <= #1 3'sb010; $display(";A 423");		//(= P1_P1_P1_State    0b010)) ;423
                        end
                        else begin
                            $display(";A 422");		//(= (bv-and (bv-comp P1_P1_P1_HOLD  0b0) (bv-comp P1_P1_P1_RequestPending  0b1))   0b0)) ;422
                            if (((P1_P1_P1_HOLD == 1'b0) & (P1_P1_P1_RequestPending == 1'b0))) begin
                                $display(";A 424");		//(= (bv-and (bv-comp P1_P1_P1_HOLD  0b0) (bv-comp P1_P1_P1_RequestPending  0b0))   0b1)) ;424
                                P1_P1_P1_State <= #1 3'sb001; $display(";A 426");		//(= P1_P1_P1_State    0b001)) ;426
                            end
                            else begin
                                $display(";A 425");		//(= (bv-and (bv-comp P1_P1_P1_HOLD  0b0) (bv-comp P1_P1_P1_RequestPending  0b0))   0b0)) ;425
                                P1_P1_P1_State <= #1 3'sb101; $display(";A 427");		//(= P1_P1_P1_State    0b101)) ;427
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 428");		//(= P1_P1_P1_State    0b110)) ;428
                        P1_P1_P1_Address <= #1 ((P1_P1_P1_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 429");		//(= P1_P1_P1_Address    (bv-smod (bv-sdiv P1_P1_P1_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;429
                        P1_P1_P1_BE_n <= #1 P1_P1_P1_ByteEnable; $display(";A 430");		//(= P1_P1_P1_BE_n    P1_P1_P1_ByteEnable )) ;430
                        P1_P1_P1_M_IO_n <= #1 P1_P1_P1_MemoryFetch; $display(";A 431");		//(= P1_P1_P1_M_IO_n    P1_P1_P1_MemoryFetch )) ;431
                        if ((P1_P1_P1_ReadRequest == 1'b1)) begin
                            $display(";A 432");		//(= (bv-comp P1_P1_P1_ReadRequest  0b1)   0b1)) ;432
                            P1_P1_P1_W_R_n <= #1 1'b0; $display(";A 434");		//(= P1_P1_P1_W_R_n    0b0)) ;434
                        end
                        else begin
                            $display(";A 433");		//(= (bv-comp P1_P1_P1_ReadRequest  0b1)   0b0)) ;433
                            P1_P1_P1_W_R_n <= #1 1'b1; $display(";A 435");		//(= P1_P1_P1_W_R_n    0b1)) ;435
                        end
                        if ((P1_P1_P1_CodeFetch == 1'b1)) begin
                            $display(";A 436");		//(= (bv-comp P1_P1_P1_CodeFetch  0b1)   0b1)) ;436
                            P1_P1_P1_D_C_n <= #1 1'b0; $display(";A 438");		//(= P1_P1_P1_D_C_n    0b0)) ;438
                        end
                        else begin
                            $display(";A 437");		//(= (bv-comp P1_P1_P1_CodeFetch  0b1)   0b0)) ;437
                            P1_P1_P1_D_C_n <= #1 1'b1; $display(";A 439");		//(= P1_P1_P1_D_C_n    0b1)) ;439
                        end
                        P1_P1_P1_ADS_n <= #1 1'b0; $display(";A 440");		//(= P1_P1_P1_ADS_n    0b0)) ;440
                        if ((P1_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 441");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;441
                            P1_P1_P1_State <= #1 3'sb100; $display(";A 443");		//(= P1_P1_P1_State    0b100)) ;443
                        end
                        else begin
                            $display(";A 442");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;442
                            P1_P1_P1_State <= #1 3'sb110; $display(";A 444");		//(= P1_P1_P1_State    0b110)) ;444
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 445");		//(= P1_P1_P1_State    0b111)) ;445
                        if ((((P1_P1_P1_READY_n == 1'b1) & (P1_P1_P1_RequestPending == 1'b1)) & (P1_P1_P1_HOLD == 1'b0))) begin
                            $display(";A 446");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b1) (bv-comp P1_P1_P1_RequestPending  0b1)) (bv-comp P1_P1_P1_HOLD  0b0))   0b1)) ;446
                            P1_P1_P1_State <= #1 3'sb110; $display(";A 448");		//(= P1_P1_P1_State    0b110)) ;448
                        end
                        else begin
                            $display(";A 447");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b1) (bv-comp P1_P1_P1_RequestPending  0b1)) (bv-comp P1_P1_P1_HOLD  0b0))   0b0)) ;447
                            if (((P1_P1_P1_READY_n == 1'b0) & (P1_P1_P1_HOLD == 1'b1))) begin
                                $display(";A 449");		//(= (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b1))   0b1)) ;449
                                P1_P1_P1_State <= #1 3'sb101; $display(";A 451");		//(= P1_P1_P1_State    0b101)) ;451
                            end
                            else begin
                                $display(";A 450");		//(= (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b1))   0b0)) ;450
                                if ((((P1_P1_P1_READY_n == 1'b0) & (P1_P1_P1_HOLD == 1'b0)) & (P1_P1_P1_RequestPending == 1'b1))) begin
                                    $display(";A 452");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b1))   0b1)) ;452
                                    P1_P1_P1_State <= #1 3'sb010; $display(";A 454");		//(= P1_P1_P1_State    0b010)) ;454
                                end
                                else begin
                                    $display(";A 453");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b1))   0b0)) ;453
                                    if ((((P1_P1_P1_READY_n == 1'b0) & (P1_P1_P1_HOLD == 1'b0)) & (P1_P1_P1_RequestPending == 1'b0))) begin
                                        $display(";A 455");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b0))   0b1)) ;455
                                        P1_P1_P1_State <= #1 3'sb001; $display(";A 457");		//(= P1_P1_P1_State    0b001)) ;457
                                    end
                                    else begin
                                        $display(";A 456");		//(= (bv-and (bv-and (bv-comp P1_P1_P1_READY_n  0b0) (bv-comp P1_P1_P1_HOLD  0b0)) (bv-comp P1_P1_P1_RequestPending  0b0))   0b0)) ;456
                                        P1_P1_P1_State <= #1 3'sb111; $display(";A 458");		//(= P1_P1_P1_State    0b111)) ;458
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:488
    always @(posedge P1_P1_P1_RESET or posedge P1_P1_P1_CLOCK) begin
        if ((P1_P1_P1_RESET == 1'b1)) begin
            $display(";A 459");		//(= (bv-comp P1_P1_P1_RESET  0b1)   0b1)) ;459
            P1_P1_P1_State2 = 4'sb0000; $display(";A 461");		//(= P1_P1_P1_State2    0b0000)) ;461
            P1_P1_P1_InstQueue[0] = 8'b00000000; $display(";A 462");		//(= P1_P1_P1_InstQueue    0b00000000)) ;462
            P1_P1_P1_InstQueue[1] = 8'b00000000; $display(";A 463");		//(= P1_P1_P1_InstQueue    0b00000000)) ;463
            P1_P1_P1_InstQueue[2] = 8'b00000000; $display(";A 464");		//(= P1_P1_P1_InstQueue    0b00000000)) ;464
            P1_P1_P1_InstQueue[3] = 8'b00000000; $display(";A 465");		//(= P1_P1_P1_InstQueue    0b00000000)) ;465
            P1_P1_P1_InstQueue[4] = 8'b00000000; $display(";A 466");		//(= P1_P1_P1_InstQueue    0b00000000)) ;466
            P1_P1_P1_InstQueue[5] = 8'b00000000; $display(";A 467");		//(= P1_P1_P1_InstQueue    0b00000000)) ;467
            P1_P1_P1_InstQueue[6] = 8'b00000000; $display(";A 468");		//(= P1_P1_P1_InstQueue    0b00000000)) ;468
            P1_P1_P1_InstQueue[7] = 8'b00000000; $display(";A 469");		//(= P1_P1_P1_InstQueue    0b00000000)) ;469
            P1_P1_P1_InstQueue[8] = 8'b00000000; $display(";A 470");		//(= P1_P1_P1_InstQueue    0b00000000)) ;470
            P1_P1_P1_InstQueue[9] = 8'b00000000; $display(";A 471");		//(= P1_P1_P1_InstQueue    0b00000000)) ;471
            P1_P1_P1_InstQueue[10] = 8'b00000000; $display(";A 472");		//(= P1_P1_P1_InstQueue    0b00000000)) ;472
            P1_P1_P1_InstQueue[11] = 8'b00000000; $display(";A 473");		//(= P1_P1_P1_InstQueue    0b00000000)) ;473
            P1_P1_P1_InstQueue[12] = 8'b00000000; $display(";A 474");		//(= P1_P1_P1_InstQueue    0b00000000)) ;474
            P1_P1_P1_InstQueue[13] = 8'b00000000; $display(";A 475");		//(= P1_P1_P1_InstQueue    0b00000000)) ;475
            P1_P1_P1_InstQueue[14] = 8'b00000000; $display(";A 476");		//(= P1_P1_P1_InstQueue    0b00000000)) ;476
            P1_P1_P1_InstQueue[15] = 8'b00000000; $display(";A 477");		//(= P1_P1_P1_InstQueue    0b00000000)) ;477
            P1_P1_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 478");		//(= P1_P1_P1_InstQueueRd_Addr    0b00000)) ;478
            P1_P1_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 479");		//(= P1_P1_P1_InstQueueWr_Addr    0b00000)) ;479
            P1_P1_P1_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 480");		//(= P1_P1_P1_InstAddrPointer    0b00000000000000000000000000000000)) ;480
            P1_P1_P1_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 481");		//(= P1_P1_P1_PhyAddrPointer    0b00000000000000000000000000000000)) ;481
            P1_P1_P1_Extended = 1'b0; $display(";A 482");		//(= P1_P1_P1_Extended    0b0)) ;482
            P1_P1_P1_More = 1'b0; $display(";A 483");		//(= P1_P1_P1_More    0b0)) ;483
            P1_P1_P1_Flush = 1'b0; $display(";A 484");		//(= P1_P1_P1_Flush    0b0)) ;484
            P1_P1_P1_lWord = 16'sb0000000000000000; $display(";A 485");		//(= P1_P1_P1_lWord    0b0000000000000000)) ;485
            P1_P1_P1_uWord = 15'sb000000000000000; $display(";A 486");		//(= P1_P1_P1_uWord    0b000000000000000)) ;486
            P1_P1_P1_fWord = 32'sb00000000000000000000000000000000; $display(";A 487");		//(= P1_P1_P1_fWord    0b00000000000000000000000000000000)) ;487
            P1_P1_P1_CodeFetch <= #1 1'b0; $display(";A 488");		//(= P1_P1_P1_CodeFetch    0b0)) ;488
            P1_P1_P1_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 489");		//(= P1_P1_P1_Datao    0b00000000000000000000000000000000)) ;489
            P1_P1_P1_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 490");		//(= P1_P1_P1_EAX    0b00000000000000000000000000000000)) ;490
            P1_P1_P1_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 491");		//(= P1_P1_P1_EBX    0b00000000000000000000000000000000)) ;491
            P1_P1_P1_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 492");		//(= P1_P1_P1_rEIP    0b00000000000000000000000000000000)) ;492
            P1_P1_P1_ReadRequest <= #1 1'b0; $display(";A 493");		//(= P1_P1_P1_ReadRequest    0b0)) ;493
            P1_P1_P1_MemoryFetch <= #1 1'b0; $display(";A 494");		//(= P1_P1_P1_MemoryFetch    0b0)) ;494
            P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 495");		//(= P1_P1_P1_RequestPending    0b0)) ;495
        end
        else begin
            $display(";A 460");		//(= (bv-comp P1_P1_P1_RESET  0b1)   0b0)) ;460
            case (P1_P1_P1_State2)
                4'b0000 :
                    begin
                        $display(";A 496");		//(= P1_P1_P1_State2    0b0000)) ;496
                        P1_P1_P1_PhyAddrPointer = P1_P1_P1_rEIP; $display(";A 497");		//(= P1_P1_P1_PhyAddrPointer    P1_P1_P1_rEIP )) ;497
                        P1_P1_P1_InstAddrPointer = P1_P1_P1_PhyAddrPointer; $display(";A 498");		//(= P1_P1_P1_InstAddrPointer    P1_P1_P1_PhyAddrPointer )) ;498
                        P1_P1_P1_State2 = 4'sb0001; $display(";A 499");		//(= P1_P1_P1_State2    0b0001)) ;499
                        P1_P1_P1_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 500");		//(= P1_P1_P1_rEIP    0b00000000000011111111111111110000)) ;500
                        P1_P1_P1_ReadRequest <= #1 1'b1; $display(";A 501");		//(= P1_P1_P1_ReadRequest    0b1)) ;501
                        P1_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 502");		//(= P1_P1_P1_MemoryFetch    0b1)) ;502
                        P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 503");		//(= P1_P1_P1_RequestPending    0b1)) ;503
                    end
                4'b0001 :
                    begin
                        $display(";A 504");		//(= P1_P1_P1_State2    0b0001)) ;504
                        P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 505");		//(= P1_P1_P1_RequestPending    0b1)) ;505
                        P1_P1_P1_ReadRequest <= #1 1'b1; $display(";A 506");		//(= P1_P1_P1_ReadRequest    0b1)) ;506
                        P1_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 507");		//(= P1_P1_P1_MemoryFetch    0b1)) ;507
                        P1_P1_P1_CodeFetch <= #1 1'b1; $display(";A 508");		//(= P1_P1_P1_CodeFetch    0b1)) ;508
                        if ((P1_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 509");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;509
                            P1_P1_P1_State2 = 4'sb0010; $display(";A 511");		//(= P1_P1_P1_State2    0b0010)) ;511
                        end
                        else begin
                            $display(";A 510");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;510
                            P1_P1_P1_State2 = 4'sb0001; $display(";A 512");		//(= P1_P1_P1_State2    0b0001)) ;512
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 513");		//(= P1_P1_P1_State2    0b0010)) ;513
                        P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 514");		//(= P1_P1_P1_RequestPending    0b0)) ;514
                        P1_P1_P1_InstQueue[P1_P1_P1_InstQueueWr_Addr] = (P1_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 515");		//(= P1_P1_P1_InstQueue    (bv-smod P1_P1_P1_Datai  0b00000000000000000000000100000000))) ;515
                        P1_P1_P1_InstQueueWr_Addr = ((P1_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 516");		//(= P1_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;516
                        P1_P1_P1_InstQueue[P1_P1_P1_InstQueueWr_Addr] = (P1_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 517");		//(= P1_P1_P1_InstQueue    (bv-smod P1_P1_P1_Datai  0b00000000000000000000000100000000))) ;517
                        P1_P1_P1_InstQueueWr_Addr = ((P1_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 518");		//(= P1_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;518
                        if ((P1_P1_P1_StateBS16 == 1'b1)) begin
                            $display(";A 519");		//(= (bv-comp P1_P1_P1_StateBS16  0b1)   0b1)) ;519
                            P1_P1_P1_InstQueue[P1_P1_P1_InstQueueWr_Addr] = ((P1_P1_P1_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 521");		//(= P1_P1_P1_InstQueue    (bv-smod (bv-sdiv P1_P1_P1_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;521
                            P1_P1_P1_InstQueueWr_Addr = ((P1_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 522");		//(= P1_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;522
                            P1_P1_P1_InstQueue[P1_P1_P1_InstQueueWr_Addr] = ((P1_P1_P1_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 523");		//(= P1_P1_P1_InstQueue    (bv-smod (bv-sdiv P1_P1_P1_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;523
                            P1_P1_P1_InstQueueWr_Addr = ((P1_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 524");		//(= P1_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;524
                            P1_P1_P1_PhyAddrPointer = (P1_P1_P1_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 525");		//(= P1_P1_P1_PhyAddrPointer    (bv-add P1_P1_P1_PhyAddrPointer  0b00000000000000000000000000000100))) ;525
                            P1_P1_P1_State2 = 4'sb0101; $display(";A 526");		//(= P1_P1_P1_State2    0b0101)) ;526
                        end
                        else begin
                            $display(";A 520");		//(= (bv-comp P1_P1_P1_StateBS16  0b1)   0b0)) ;520
                            P1_P1_P1_PhyAddrPointer = (P1_P1_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 527");		//(= P1_P1_P1_PhyAddrPointer    (bv-add P1_P1_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;527
                            if ((P1_P1_P1_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 528");		//(= (bool-to-bv (bv-slt P1_P1_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;528
                                P1_P1_P1_rEIP <= #1 (-P1_P1_P1_PhyAddrPointer); $display(";A 530");		//(= P1_P1_P1_rEIP    (bv-neg P1_P1_P1_PhyAddrPointer ))) ;530
                            end
                            else begin
                                $display(";A 529");		//(= (bool-to-bv (bv-slt P1_P1_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;529
                                P1_P1_P1_rEIP <= #1 P1_P1_P1_PhyAddrPointer; $display(";A 531");		//(= P1_P1_P1_rEIP    P1_P1_P1_PhyAddrPointer )) ;531
                            end
                            P1_P1_P1_State2 = 4'sb0011; $display(";A 532");		//(= P1_P1_P1_State2    0b0011)) ;532
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 533");		//(= P1_P1_P1_State2    0b0011)) ;533
                        P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 534");		//(= P1_P1_P1_RequestPending    0b1)) ;534
                        if ((P1_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 535");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;535
                            P1_P1_P1_State2 = 4'sb0100; $display(";A 537");		//(= P1_P1_P1_State2    0b0100)) ;537
                        end
                        else begin
                            $display(";A 536");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;536
                            P1_P1_P1_State2 = 4'sb0011; $display(";A 538");		//(= P1_P1_P1_State2    0b0011)) ;538
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 539");		//(= P1_P1_P1_State2    0b0100)) ;539
                        P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 540");		//(= P1_P1_P1_RequestPending    0b0)) ;540
                        P1_P1_P1_InstQueue[P1_P1_P1_InstQueueWr_Addr] = (P1_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 541");		//(= P1_P1_P1_InstQueue    (bv-smod P1_P1_P1_Datai  0b00000000000000000000000100000000))) ;541
                        P1_P1_P1_InstQueueWr_Addr = ((P1_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 542");		//(= P1_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;542
                        P1_P1_P1_InstQueue[P1_P1_P1_InstQueueWr_Addr] = (P1_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 543");		//(= P1_P1_P1_InstQueue    (bv-smod P1_P1_P1_Datai  0b00000000000000000000000100000000))) ;543
                        P1_P1_P1_InstQueueWr_Addr = ((P1_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 544");		//(= P1_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;544
                        P1_P1_P1_PhyAddrPointer = (P1_P1_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 545");		//(= P1_P1_P1_PhyAddrPointer    (bv-add P1_P1_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;545
                        P1_P1_P1_State2 = 4'sb0101; $display(";A 546");		//(= P1_P1_P1_State2    0b0101)) ;546
                    end
                4'b0101 :
                    begin
                        $display(";A 547");		//(= P1_P1_P1_State2    0b0101)) ;547
                        case (P1_P1_P1_InstQueue[P1_P1_P1_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 548");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b10010000)) ;548
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 549");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;549
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 550");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;550
                                    P1_P1_P1_Flush = 1'b0; $display(";A 551");		//(= P1_P1_P1_Flush    0b0)) ;551
                                    P1_P1_P1_More = 1'b0; $display(";A 552");		//(= P1_P1_P1_More    0b0)) ;552
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 553");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b01100110)) ;553
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 554");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;554
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 555");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;555
                                    P1_P1_P1_Extended = 1'b1; $display(";A 556");		//(= P1_P1_P1_Extended    0b1)) ;556
                                    P1_P1_P1_Flush = 1'b0; $display(";A 557");		//(= P1_P1_P1_Flush    0b0)) ;557
                                    P1_P1_P1_More = 1'b0; $display(";A 558");		//(= P1_P1_P1_More    0b0)) ;558
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 559");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b11101011)) ;559
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 560");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;560
                                        if ((P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 562");		//(= (bool-to-bv (bv-gt P1_P1_P1_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;562
                                            P1_P1_P1_PhyAddrPointer = ((P1_P1_P1_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 564");		//(= P1_P1_P1_PhyAddrPointer    (bv-sub (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P1_P1_P1_InstQueue 0 )))) ;564
                                            P1_P1_P1_InstAddrPointer = P1_P1_P1_PhyAddrPointer; $display(";A 565");		//(= P1_P1_P1_InstAddrPointer    P1_P1_P1_PhyAddrPointer )) ;565
                                        end
                                        else begin
                                            $display(";A 563");		//(= (bool-to-bv (bv-gt P1_P1_P1_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;563
                                            P1_P1_P1_PhyAddrPointer = ((P1_P1_P1_InstAddrPointer + 32'b00000000000000000000000000000010) + P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 566");		//(= P1_P1_P1_PhyAddrPointer    (bv-add (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000010) P1_P1_P1_InstQueue 0 ))) ;566
                                            P1_P1_P1_InstAddrPointer = P1_P1_P1_PhyAddrPointer; $display(";A 567");		//(= P1_P1_P1_InstAddrPointer    P1_P1_P1_PhyAddrPointer )) ;567
                                        end
                                        P1_P1_P1_Flush = 1'b1; $display(";A 568");		//(= P1_P1_P1_Flush    0b1)) ;568
                                        P1_P1_P1_More = 1'b0; $display(";A 569");		//(= P1_P1_P1_More    0b0)) ;569
                                    end
                                    else begin
                                        $display(";A 561");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;561
                                        P1_P1_P1_Flush = 1'b0; $display(";A 570");		//(= P1_P1_P1_Flush    0b0)) ;570
                                        P1_P1_P1_More = 1'b1; $display(";A 571");		//(= P1_P1_P1_More    0b1)) ;571
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 572");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b11101001)) ;572
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 573");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;573
                                        P1_P1_P1_PhyAddrPointer = ((P1_P1_P1_InstAddrPointer + 32'b00000000000000000000000000000101) + P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 575");		//(= P1_P1_P1_PhyAddrPointer    (bv-add (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000101) P1_P1_P1_InstQueue 0 ))) ;575
                                        P1_P1_P1_InstAddrPointer = P1_P1_P1_PhyAddrPointer; $display(";A 576");		//(= P1_P1_P1_InstAddrPointer    P1_P1_P1_PhyAddrPointer )) ;576
                                        P1_P1_P1_Flush = 1'b1; $display(";A 577");		//(= P1_P1_P1_Flush    0b1)) ;577
                                        P1_P1_P1_More = 1'b0; $display(";A 578");		//(= P1_P1_P1_More    0b0)) ;578
                                    end
                                    else begin
                                        $display(";A 574");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;574
                                        P1_P1_P1_Flush = 1'b0; $display(";A 579");		//(= P1_P1_P1_Flush    0b0)) ;579
                                        P1_P1_P1_More = 1'b1; $display(";A 580");		//(= P1_P1_P1_More    0b1)) ;580
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 581");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b11101010)) ;581
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 582");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;582
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 583");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;583
                                    P1_P1_P1_Flush = 1'b0; $display(";A 584");		//(= P1_P1_P1_Flush    0b0)) ;584
                                    P1_P1_P1_More = 1'b0; $display(";A 585");		//(= P1_P1_P1_More    0b0)) ;585
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 586");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b10110000)) ;586
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 587");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;587
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 588");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;588
                                    P1_P1_P1_Flush = 1'b0; $display(";A 589");		//(= P1_P1_P1_Flush    0b0)) ;589
                                    P1_P1_P1_More = 1'b0; $display(";A 590");		//(= P1_P1_P1_More    0b0)) ;590
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 591");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b10111000)) ;591
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 592");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;592
                                        P1_P1_P1_EAX <= #1 ((((P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 594");		//(= P1_P1_P1_EAX    (bv-add (bv-add (bv-add (bv-mul P1_P1_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P1_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P1_P1_InstQueue 0  0b00000000000000000000000100000000)) P1_P1_P1_InstQueue 0 ))) ;594
                                        P1_P1_P1_More = 1'b0; $display(";A 595");		//(= P1_P1_P1_More    0b0)) ;595
                                        P1_P1_P1_Flush = 1'b0; $display(";A 596");		//(= P1_P1_P1_Flush    0b0)) ;596
                                        P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 597");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;597
                                        P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 598");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;598
                                    end
                                    else begin
                                        $display(";A 593");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;593
                                        P1_P1_P1_Flush = 1'b0; $display(";A 599");		//(= P1_P1_P1_Flush    0b0)) ;599
                                        P1_P1_P1_More = 1'b1; $display(";A 600");		//(= P1_P1_P1_More    0b1)) ;600
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 601");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b10111011)) ;601
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 602");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;602
                                        P1_P1_P1_EBX <= #1 ((((P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P1_P1_InstQueue[((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 604");		//(= P1_P1_P1_EBX    (bv-add (bv-add (bv-add (bv-mul P1_P1_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P1_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P1_P1_InstQueue 0  0b00000000000000000000000100000000)) P1_P1_P1_InstQueue 0 ))) ;604
                                        P1_P1_P1_More = 1'b0; $display(";A 605");		//(= P1_P1_P1_More    0b0)) ;605
                                        P1_P1_P1_Flush = 1'b0; $display(";A 606");		//(= P1_P1_P1_Flush    0b0)) ;606
                                        P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 607");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;607
                                        P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 608");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;608
                                    end
                                    else begin
                                        $display(";A 603");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;603
                                        P1_P1_P1_Flush = 1'b0; $display(";A 609");		//(= P1_P1_P1_Flush    0b0)) ;609
                                        P1_P1_P1_More = 1'b1; $display(";A 610");		//(= P1_P1_P1_More    0b1)) ;610
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 611");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b10001011)) ;611
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 612");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;612
                                        if ((P1_P1_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 614");		//(= (bool-to-bv (bv-slt P1_P1_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;614
                                            P1_P1_P1_rEIP <= #1 (-P1_P1_P1_EBX); $display(";A 616");		//(= P1_P1_P1_rEIP    (bv-neg P1_P1_P1_EBX ))) ;616
                                        end
                                        else begin
                                            $display(";A 615");		//(= (bool-to-bv (bv-slt P1_P1_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;615
                                            P1_P1_P1_rEIP <= #1 P1_P1_P1_EBX; $display(";A 617");		//(= P1_P1_P1_rEIP    P1_P1_P1_EBX )) ;617
                                        end
                                        P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 618");		//(= P1_P1_P1_RequestPending    0b1)) ;618
                                        P1_P1_P1_ReadRequest <= #1 1'b1; $display(";A 619");		//(= P1_P1_P1_ReadRequest    0b1)) ;619
                                        P1_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 620");		//(= P1_P1_P1_MemoryFetch    0b1)) ;620
                                        P1_P1_P1_CodeFetch <= #1 1'b0; $display(";A 621");		//(= P1_P1_P1_CodeFetch    0b0)) ;621
                                        if ((P1_P1_P1_READY_n == 1'b0)) begin
                                            $display(";A 622");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;622
                                            P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 624");		//(= P1_P1_P1_RequestPending    0b0)) ;624
                                            P1_P1_P1_uWord = (P1_P1_P1_Datai % 32'b00000000000000001000000000000000); $display(";A 625");		//(= P1_P1_P1_uWord    (bv-smod P1_P1_P1_Datai  0b00000000000000001000000000000000))) ;625
                                            if ((P1_P1_P1_StateBS16 == 1'b1)) begin
                                                $display(";A 626");		//(= (bv-comp P1_P1_P1_StateBS16  0b1)   0b1)) ;626
                                                P1_P1_P1_lWord = (P1_P1_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 628");		//(= P1_P1_P1_lWord    (bv-smod P1_P1_P1_Datai  0b00000000000000010000000000000000))) ;628
                                            end
                                            else begin
                                                $display(";A 627");		//(= (bv-comp P1_P1_P1_StateBS16  0b1)   0b0)) ;627
                                                P1_P1_P1_rEIP <= #1 (P1_P1_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 629");		//(= P1_P1_P1_rEIP    (bv-add P1_P1_P1_rEIP  0b00000000000000000000000000000010))) ;629
                                                P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 630");		//(= P1_P1_P1_RequestPending    0b1)) ;630
                                                if ((P1_P1_P1_READY_n == 1'b0)) begin
                                                    $display(";A 631");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;631
                                                    P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 633");		//(= P1_P1_P1_RequestPending    0b0)) ;633
                                                    P1_P1_P1_lWord = (P1_P1_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 634");		//(= P1_P1_P1_lWord    (bv-smod P1_P1_P1_Datai  0b00000000000000010000000000000000))) ;634
                                                end
                                                else begin
                                                    $display(";A 632");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;632
                                                end
                                            end
                                            if ((P1_P1_P1_READY_n == 1'b0)) begin
                                                $display(";A 635");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;635
                                                P1_P1_P1_EAX <= #1 ((P1_P1_P1_uWord * 32'b00000000000000010000000000000000) + P1_P1_P1_lWord); $display(";A 637");		//(= P1_P1_P1_EAX    (bv-add (bv-mul P1_P1_P1_uWord  0b00000000000000010000000000000000) P1_P1_P1_lWord ))) ;637
                                                P1_P1_P1_More = 1'b0; $display(";A 638");		//(= P1_P1_P1_More    0b0)) ;638
                                                P1_P1_P1_Flush = 1'b0; $display(";A 639");		//(= P1_P1_P1_Flush    0b0)) ;639
                                                P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 640");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;640
                                                P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 641");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;641
                                            end
                                            else begin
                                                $display(";A 636");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;636
                                            end
                                        end
                                        else begin
                                            $display(";A 623");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;623
                                        end
                                    end
                                    else begin
                                        $display(";A 613");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;613
                                        P1_P1_P1_Flush = 1'b0; $display(";A 642");		//(= P1_P1_P1_Flush    0b0)) ;642
                                        P1_P1_P1_More = 1'b1; $display(";A 643");		//(= P1_P1_P1_More    0b1)) ;643
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 644");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b10001001)) ;644
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 645");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;645
                                        if ((P1_P1_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 647");		//(= (bool-to-bv (bv-slt P1_P1_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;647
                                            P1_P1_P1_rEIP <= #1 P1_P1_P1_EBX; $display(";A 649");		//(= P1_P1_P1_rEIP    P1_P1_P1_EBX )) ;649
                                        end
                                        else begin
                                            $display(";A 648");		//(= (bool-to-bv (bv-slt P1_P1_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;648
                                            P1_P1_P1_rEIP <= #1 P1_P1_P1_EBX; $display(";A 650");		//(= P1_P1_P1_rEIP    P1_P1_P1_EBX )) ;650
                                        end
                                        P1_P1_P1_lWord = (P1_P1_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 651");		//(= P1_P1_P1_lWord    (bv-smod P1_P1_P1_EAX  0b00000000000000010000000000000000))) ;651
                                        P1_P1_P1_uWord = ((P1_P1_P1_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 652");		//(= P1_P1_P1_uWord    (bv-smod (bv-sdiv P1_P1_P1_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;652
                                        P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 653");		//(= P1_P1_P1_RequestPending    0b1)) ;653
                                        P1_P1_P1_ReadRequest <= #1 1'b0; $display(";A 654");		//(= P1_P1_P1_ReadRequest    0b0)) ;654
                                        P1_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 655");		//(= P1_P1_P1_MemoryFetch    0b1)) ;655
                                        P1_P1_P1_CodeFetch <= #1 1'b0; $display(";A 656");		//(= P1_P1_P1_CodeFetch    0b0)) ;656
                                        if (((P1_P1_P1_State == 32'b00000000000000000000000000000010) | (P1_P1_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 657");		//(= (bv-or (bv-comp P1_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P1_State  0b00000000000000000000000000000100))   0b1)) ;657
                                            P1_P1_P1_Datao <= #1 ((P1_P1_P1_uWord * 32'b00000000000000010000000000000000) + P1_P1_P1_lWord); $display(";A 659");		//(= P1_P1_P1_Datao    (bv-add (bv-mul P1_P1_P1_uWord  0b00000000000000010000000000000000) P1_P1_P1_lWord ))) ;659
                                            if ((P1_P1_P1_READY_n == 1'b0)) begin
                                                $display(";A 660");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;660
                                                P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 662");		//(= P1_P1_P1_RequestPending    0b0)) ;662
                                                if ((P1_P1_P1_StateBS16 == 1'b0)) begin
                                                    $display(";A 663");		//(= (bv-comp P1_P1_P1_StateBS16  0b0)   0b1)) ;663
                                                    P1_P1_P1_rEIP <= #1 (P1_P1_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 665");		//(= P1_P1_P1_rEIP    (bv-add P1_P1_P1_rEIP  0b00000000000000000000000000000010))) ;665
                                                    P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 666");		//(= P1_P1_P1_RequestPending    0b1)) ;666
                                                    P1_P1_P1_ReadRequest <= #1 1'b0; $display(";A 667");		//(= P1_P1_P1_ReadRequest    0b0)) ;667
                                                    P1_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 668");		//(= P1_P1_P1_MemoryFetch    0b1)) ;668
                                                    P1_P1_P1_CodeFetch <= #1 1'b0; $display(";A 669");		//(= P1_P1_P1_CodeFetch    0b0)) ;669
                                                    P1_P1_P1_State2 = 4'sb0110; $display(";A 670");		//(= P1_P1_P1_State2    0b0110)) ;670
                                                end
                                                else begin
                                                    $display(";A 664");		//(= (bv-comp P1_P1_P1_StateBS16  0b0)   0b0)) ;664
                                                end
                                                P1_P1_P1_More = 1'b0; $display(";A 671");		//(= P1_P1_P1_More    0b0)) ;671
                                                P1_P1_P1_Flush = 1'b0; $display(";A 672");		//(= P1_P1_P1_Flush    0b0)) ;672
                                                P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 673");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;673
                                                P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 674");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;674
                                            end
                                            else begin
                                                $display(";A 661");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;661
                                            end
                                        end
                                        else begin
                                            $display(";A 658");		//(= (bv-or (bv-comp P1_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P1_State  0b00000000000000000000000000000100))   0b0)) ;658
                                        end
                                    end
                                    else begin
                                        $display(";A 646");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;646
                                        P1_P1_P1_Flush = 1'b0; $display(";A 675");		//(= P1_P1_P1_Flush    0b0)) ;675
                                        P1_P1_P1_More = 1'b1; $display(";A 676");		//(= P1_P1_P1_More    0b1)) ;676
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 677");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b11100100)) ;677
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 678");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;678
                                        P1_P1_P1_rEIP <= #1 (P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 680");		//(= P1_P1_P1_rEIP    (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;680
                                        P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 681");		//(= P1_P1_P1_RequestPending    0b1)) ;681
                                        P1_P1_P1_ReadRequest <= #1 1'b1; $display(";A 682");		//(= P1_P1_P1_ReadRequest    0b1)) ;682
                                        P1_P1_P1_MemoryFetch <= #1 1'b0; $display(";A 683");		//(= P1_P1_P1_MemoryFetch    0b0)) ;683
                                        P1_P1_P1_CodeFetch <= #1 1'b0; $display(";A 684");		//(= P1_P1_P1_CodeFetch    0b0)) ;684
                                        if ((P1_P1_P1_READY_n == 1'b0)) begin
                                            $display(";A 685");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;685
                                            P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 687");		//(= P1_P1_P1_RequestPending    0b0)) ;687
                                            P1_P1_P1_EAX <= #1 P1_P1_P1_Datai; $display(";A 688");		//(= P1_P1_P1_EAX    P1_P1_P1_Datai )) ;688
                                            P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 689");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;689
                                            P1_P1_P1_InstQueueRd_Addr = (P1_P1_P1_InstQueueRd_Addr + 5'b00010); $display(";A 690");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-add P1_P1_P1_InstQueueRd_Addr  0b00010))) ;690
                                            P1_P1_P1_Flush = 1'b0; $display(";A 691");		//(= P1_P1_P1_Flush    0b0)) ;691
                                            P1_P1_P1_More = 1'b0; $display(";A 692");		//(= P1_P1_P1_More    0b0)) ;692
                                        end
                                        else begin
                                            $display(";A 686");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;686
                                        end
                                    end
                                    else begin
                                        $display(";A 679");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;679
                                        P1_P1_P1_Flush = 1'b0; $display(";A 693");		//(= P1_P1_P1_Flush    0b0)) ;693
                                        P1_P1_P1_More = 1'b1; $display(";A 694");		//(= P1_P1_P1_More    0b1)) ;694
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 695");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b11100110)) ;695
                                    if (((P1_P1_P1_InstQueueWr_Addr - P1_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 696");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;696
                                        P1_P1_P1_rEIP <= #1 (P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 698");		//(= P1_P1_P1_rEIP    (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;698
                                        P1_P1_P1_RequestPending <= #1 1'b1; $display(";A 699");		//(= P1_P1_P1_RequestPending    0b1)) ;699
                                        P1_P1_P1_ReadRequest <= #1 1'b0; $display(";A 700");		//(= P1_P1_P1_ReadRequest    0b0)) ;700
                                        P1_P1_P1_MemoryFetch <= #1 1'b0; $display(";A 701");		//(= P1_P1_P1_MemoryFetch    0b0)) ;701
                                        P1_P1_P1_CodeFetch <= #1 1'b0; $display(";A 702");		//(= P1_P1_P1_CodeFetch    0b0)) ;702
                                        if (((P1_P1_P1_State == 32'b00000000000000000000000000000010) | (P1_P1_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 703");		//(= (bv-or (bv-comp P1_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P1_State  0b00000000000000000000000000000100))   0b1)) ;703
                                            P1_P1_P1_fWord = (P1_P1_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 705");		//(= P1_P1_P1_fWord    (bv-smod P1_P1_P1_EAX  0b00000000000000010000000000000000))) ;705
                                            P1_P1_P1_Datao <= #1 P1_P1_P1_fWord; $display(";A 706");		//(= P1_P1_P1_Datao    P1_P1_P1_fWord )) ;706
                                            if ((P1_P1_P1_READY_n == 1'b0)) begin
                                                $display(";A 707");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;707
                                                P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 709");		//(= P1_P1_P1_RequestPending    0b0)) ;709
                                                P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 710");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;710
                                                P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 711");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;711
                                                P1_P1_P1_Flush = 1'b0; $display(";A 712");		//(= P1_P1_P1_Flush    0b0)) ;712
                                                P1_P1_P1_More = 1'b0; $display(";A 713");		//(= P1_P1_P1_More    0b0)) ;713
                                            end
                                            else begin
                                                $display(";A 708");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;708
                                            end
                                        end
                                        else begin
                                            $display(";A 704");		//(= (bv-or (bv-comp P1_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P1_State  0b00000000000000000000000000000100))   0b0)) ;704
                                        end
                                    end
                                    else begin
                                        $display(";A 697");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P1_InstQueueWr_Addr  P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;697
                                        P1_P1_P1_Flush = 1'b0; $display(";A 714");		//(= P1_P1_P1_Flush    0b0)) ;714
                                        P1_P1_P1_More = 1'b1; $display(";A 715");		//(= P1_P1_P1_More    0b1)) ;715
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 716");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b00000100)) ;716
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 717");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;717
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 718");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;718
                                    P1_P1_P1_Flush = 1'b0; $display(";A 719");		//(= P1_P1_P1_Flush    0b0)) ;719
                                    P1_P1_P1_More = 1'b0; $display(";A 720");		//(= P1_P1_P1_More    0b0)) ;720
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 721");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b00000101)) ;721
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 722");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;722
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 723");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;723
                                    P1_P1_P1_Flush = 1'b0; $display(";A 724");		//(= P1_P1_P1_Flush    0b0)) ;724
                                    P1_P1_P1_More = 1'b0; $display(";A 725");		//(= P1_P1_P1_More    0b0)) ;725
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 726");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b11010000)) ;726
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 727");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;727
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 728");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;728
                                    P1_P1_P1_Flush = 1'b0; $display(";A 729");		//(= P1_P1_P1_Flush    0b0)) ;729
                                    P1_P1_P1_More = 1'b0; $display(";A 730");		//(= P1_P1_P1_More    0b0)) ;730
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 731");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b11000000)) ;731
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 732");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;732
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 733");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;733
                                    P1_P1_P1_Flush = 1'b0; $display(";A 734");		//(= P1_P1_P1_Flush    0b0)) ;734
                                    P1_P1_P1_More = 1'b0; $display(";A 735");		//(= P1_P1_P1_More    0b0)) ;735
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 736");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b01000000)) ;736
                                    P1_P1_P1_EAX <= #1 (P1_P1_P1_EAX + 32'sb00000000000000000000000000000001); $display(";A 737");		//(= P1_P1_P1_EAX    (bv-add P1_P1_P1_EAX  0b00000000000000000000000000000001))) ;737
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 738");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;738
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 739");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;739
                                    P1_P1_P1_Flush = 1'b0; $display(";A 740");		//(= P1_P1_P1_Flush    0b0)) ;740
                                    P1_P1_P1_More = 1'b0; $display(";A 741");		//(= P1_P1_P1_More    0b0)) ;741
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 742");		//(= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr )   0b01000011)) ;742
                                    P1_P1_P1_EBX <= #1 (P1_P1_P1_EBX + 32'sb00000000000000000000000000000001); $display(";A 743");		//(= P1_P1_P1_EBX    (bv-add P1_P1_P1_EBX  0b00000000000000000000000000000001))) ;743
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 744");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;744
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 745");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;745
                                    P1_P1_P1_Flush = 1'b0; $display(";A 746");		//(= P1_P1_P1_Flush    0b0)) ;746
                                    P1_P1_P1_More = 1'b0; $display(";A 747");		//(= P1_P1_P1_More    0b0)) ;747
                                end
                            default:
                                begin
                                    $display(";A 748");		//(= (and (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b10010000) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b01100110) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b11101011) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b11101001) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b11101010) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b10110000) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b10111000) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b10111011) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b10001011) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b10001001) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b11100100) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b11100110) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b00000100) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b00000101) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b11010000) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b11000000) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b01000000) (/= ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ) 0b01000011))   true)) ;748
                                    P1_P1_P1_InstAddrPointer = (P1_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 749");		//(= P1_P1_P1_InstAddrPointer    (bv-add P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;749
                                    P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 750");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;750
                                    P1_P1_P1_Flush = 1'b0; $display(";A 751");		//(= P1_P1_P1_Flush    0b0)) ;751
                                    P1_P1_P1_More = 1'b0; $display(";A 752");		//(= P1_P1_P1_More    0b0)) ;752
                                end
                        endcase
                        if (((~(P1_P1_P1_InstQueueRd_Addr < P1_P1_P1_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P1_P1_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P1_P1_P1_Flush) | P1_P1_P1_More))) begin
                            $display(";A 753");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P1_P1_InstQueueRd_Addr  P1_P1_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P1_P1_Flush ) P1_P1_P1_More ))   0b1)) ;753
                            P1_P1_P1_State2 = 4'sb0111; $display(";A 755");		//(= P1_P1_P1_State2    0b0111)) ;755
                        end
                        else begin
                            $display(";A 754");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P1_P1_InstQueueRd_Addr  P1_P1_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P1_P1_Flush ) P1_P1_P1_More ))   0b0)) ;754
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 756");		//(= P1_P1_P1_State2    0b0110)) ;756
                        P1_P1_P1_Datao <= #1 ((P1_P1_P1_uWord * 32'b00000000000000010000000000000000) + P1_P1_P1_lWord); $display(";A 757");		//(= P1_P1_P1_Datao    (bv-add (bv-mul P1_P1_P1_uWord  0b00000000000000010000000000000000) P1_P1_P1_lWord ))) ;757
                        if ((P1_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 758");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b1)) ;758
                            P1_P1_P1_RequestPending <= #1 1'b0; $display(";A 760");		//(= P1_P1_P1_RequestPending    0b0)) ;760
                            P1_P1_P1_State2 = 4'sb0101; $display(";A 761");		//(= P1_P1_P1_State2    0b0101)) ;761
                        end
                        else begin
                            $display(";A 759");		//(= (bv-comp P1_P1_P1_READY_n  0b0)   0b0)) ;759
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 762");		//(= P1_P1_P1_State2    0b0111)) ;762
                        if (P1_P1_P1_Flush) begin
                            $display(";A 763");		//(= P1_P1_P1_Flush    0b1)) ;763
                            P1_P1_P1_InstQueueRd_Addr = 5'sb00001; $display(";A 765");		//(= P1_P1_P1_InstQueueRd_Addr    0b00001)) ;765
                            P1_P1_P1_InstQueueWr_Addr = 5'sb00001; $display(";A 766");		//(= P1_P1_P1_InstQueueWr_Addr    0b00001)) ;766
                            if ((P1_P1_P1_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 767");		//(= (bool-to-bv (bv-slt P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;767
                                P1_P1_P1_fWord = (-P1_P1_P1_InstAddrPointer); $display(";A 769");		//(= P1_P1_P1_fWord    (bv-neg P1_P1_P1_InstAddrPointer ))) ;769
                            end
                            else begin
                                $display(";A 768");		//(= (bool-to-bv (bv-slt P1_P1_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;768
                                P1_P1_P1_fWord = P1_P1_P1_InstAddrPointer; $display(";A 770");		//(= P1_P1_P1_fWord    P1_P1_P1_InstAddrPointer )) ;770
                            end
                            if (((P1_P1_P1_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 771");		//(= (bv-comp (bv-smod P1_P1_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;771
                                P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + (P1_P1_P1_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 773");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  (bv-smod P1_P1_P1_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;773
                            end
                            else begin
                                $display(";A 772");		//(= (bv-comp (bv-smod P1_P1_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;772
                            end
                        end
                        else begin
                            $display(";A 764");		//(= P1_P1_P1_Flush    0b0)) ;764
                        end
                        if (((32'b00000000000000000000000000001111 - P1_P1_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 774");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;774
                            P1_P1_P1_State2 = 4'sb1000; $display(";A 776");		//(= P1_P1_P1_State2    0b1000)) ;776
                            P1_P1_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 777");		//(= P1_P1_P1_InstQueueWr_Addr    0b00000)) ;777
                        end
                        else begin
                            $display(";A 775");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;775
                            P1_P1_P1_State2 = 4'sb1001; $display(";A 778");		//(= P1_P1_P1_State2    0b1001)) ;778
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 779");		//(= P1_P1_P1_State2    0b1000)) ;779
                        if ((P1_P1_P1_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 780");		//(= (bool-to-bv (bv-le P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;780
                            P1_P1_P1_InstQueue[P1_P1_P1_InstQueueWr_Addr] = P1_P1_P1_InstQueue[P1_P1_P1_InstQueueRd_Addr]; $display(";A 782");		//(= P1_P1_P1_InstQueue    ( P1_P1_P1_InstQueue P1_P1_P1_InstQueueRd_Addr ))) ;782
                            P1_P1_P1_InstQueueRd_Addr = ((P1_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 783");		//(= P1_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;783
                            P1_P1_P1_InstQueueWr_Addr = ((P1_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 784");		//(= P1_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;784
                            P1_P1_P1_State2 = 4'sb1000; $display(";A 785");		//(= P1_P1_P1_State2    0b1000)) ;785
                        end
                        else begin
                            $display(";A 781");		//(= (bool-to-bv (bv-le P1_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;781
                            P1_P1_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 786");		//(= P1_P1_P1_InstQueueRd_Addr    0b00000)) ;786
                            P1_P1_P1_State2 = 4'sb1001; $display(";A 787");		//(= P1_P1_P1_State2    0b1001)) ;787
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 788");		//(= P1_P1_P1_State2    0b1001)) ;788
                        P1_P1_P1_rEIP <= #1 P1_P1_P1_PhyAddrPointer; $display(";A 789");		//(= P1_P1_P1_rEIP    P1_P1_P1_PhyAddrPointer )) ;789
                        P1_P1_P1_State2 = 4'sb0001; $display(";A 790");		//(= P1_P1_P1_State2    0b0001)) ;790
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:927
    always @(posedge P1_P1_P1_RESET or posedge P1_P1_P1_CLOCK) begin
        if ((P1_P1_P1_RESET == 1'b1)) begin
            $display(";A 791");		//(= (bv-comp P1_P1_P1_RESET  0b1)   0b1)) ;791
            P1_P1_P1_ByteEnable <= #1 4'b0000; $display(";A 793");		//(= P1_P1_P1_ByteEnable    0b0000)) ;793
            P1_P1_P1_NonAligned <= #1 1'b0; $display(";A 794");		//(= P1_P1_P1_NonAligned    0b0)) ;794
        end
        else begin
            $display(";A 792");		//(= (bv-comp P1_P1_P1_RESET  0b1)   0b0)) ;792
            case (P1_P1_P1_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 795");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000000)) ;795
                        case ((P1_P1_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 796");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;796
                                    P1_P1_P1_ByteEnable <= #1 4'b1110; $display(";A 797");		//(= P1_P1_P1_ByteEnable    0b1110)) ;797
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 798");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;798
                                    P1_P1_P1_ByteEnable <= #1 4'b1101; $display(";A 799");		//(= P1_P1_P1_ByteEnable    0b1101)) ;799
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 800");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;800
                                    P1_P1_P1_ByteEnable <= #1 4'b1011; $display(";A 801");		//(= P1_P1_P1_ByteEnable    0b1011)) ;801
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 802");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;802
                                    P1_P1_P1_ByteEnable <= #1 4'b0111; $display(";A 803");		//(= P1_P1_P1_ByteEnable    0b0111)) ;803
                                end
                            default:
                                begin
                                    $display(";A 804");		//(= (and (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;804
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 805");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000001)) ;805
                        case ((P1_P1_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 806");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;806
                                    P1_P1_P1_ByteEnable <= #1 4'b1100; $display(";A 807");		//(= P1_P1_P1_ByteEnable    0b1100)) ;807
                                    P1_P1_P1_NonAligned <= #1 1'b0; $display(";A 808");		//(= P1_P1_P1_NonAligned    0b0)) ;808
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 809");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;809
                                    P1_P1_P1_ByteEnable <= #1 4'b1001; $display(";A 810");		//(= P1_P1_P1_ByteEnable    0b1001)) ;810
                                    P1_P1_P1_NonAligned <= #1 1'b0; $display(";A 811");		//(= P1_P1_P1_NonAligned    0b0)) ;811
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 812");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;812
                                    P1_P1_P1_ByteEnable <= #1 4'b0011; $display(";A 813");		//(= P1_P1_P1_ByteEnable    0b0011)) ;813
                                    P1_P1_P1_NonAligned <= #1 1'b0; $display(";A 814");		//(= P1_P1_P1_NonAligned    0b0)) ;814
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 815");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;815
                                    P1_P1_P1_ByteEnable <= #1 4'b0111; $display(";A 816");		//(= P1_P1_P1_ByteEnable    0b0111)) ;816
                                    P1_P1_P1_NonAligned <= #1 1'b1; $display(";A 817");		//(= P1_P1_P1_NonAligned    0b1)) ;817
                                end
                            default:
                                begin
                                    $display(";A 818");		//(= (and (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;818
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 819");		//(= P1_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;819
                        case ((P1_P1_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 820");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;820
                                    P1_P1_P1_ByteEnable <= #1 4'b0000; $display(";A 821");		//(= P1_P1_P1_ByteEnable    0b0000)) ;821
                                    P1_P1_P1_NonAligned <= #1 1'b0; $display(";A 822");		//(= P1_P1_P1_NonAligned    0b0)) ;822
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 823");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;823
                                    P1_P1_P1_ByteEnable <= #1 4'b0001; $display(";A 824");		//(= P1_P1_P1_ByteEnable    0b0001)) ;824
                                    P1_P1_P1_NonAligned <= #1 1'b1; $display(";A 825");		//(= P1_P1_P1_NonAligned    0b1)) ;825
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 826");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;826
                                    P1_P1_P1_NonAligned <= #1 1'b1; $display(";A 827");		//(= P1_P1_P1_NonAligned    0b1)) ;827
                                    P1_P1_P1_ByteEnable <= #1 4'b0011; $display(";A 828");		//(= P1_P1_P1_ByteEnable    0b0011)) ;828
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 829");		//(= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;829
                                    P1_P1_P1_NonAligned <= #1 1'b1; $display(";A 830");		//(= P1_P1_P1_NonAligned    0b1)) ;830
                                    P1_P1_P1_ByteEnable <= #1 4'b0111; $display(";A 831");		//(= P1_P1_P1_ByteEnable    0b0111)) ;831
                                end
                            default:
                                begin
                                    $display(";A 832");		//(= (and (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;832
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 833");		//(= (and (/= P1_P1_P1_DataWidth  0b00000000000000000000000000000000) (/= P1_P1_P1_DataWidth  0b00000000000000000000000000000001) (/= P1_P1_P1_DataWidth  0b00000000000000000000000000000010))   true)) ;833
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:1115
    always @(posedge P1_P1_P2_RESET or posedge P1_P1_P2_CLOCK) begin
        if ((P1_P1_P2_RESET == 1'b1)) begin
            $display(";A 834");		//(= (bv-comp P1_P1_P2_RESET  0b1)   0b1)) ;834
            P1_P1_P2_BE_n <= #1 4'b0000; $display(";A 836");		//(= P1_P1_P2_BE_n    0b0000)) ;836
            P1_P1_P2_Address <= #1 30'sb000000000000000000000000000000; $display(";A 837");		//(= P1_P1_P2_Address    0b000000000000000000000000000000)) ;837
            P1_P1_P2_W_R_n <= #1 1'b0; $display(";A 838");		//(= P1_P1_P2_W_R_n    0b0)) ;838
            P1_P1_P2_D_C_n <= #1 1'b0; $display(";A 839");		//(= P1_P1_P2_D_C_n    0b0)) ;839
            P1_P1_P2_M_IO_n <= #1 1'b0; $display(";A 840");		//(= P1_P1_P2_M_IO_n    0b0)) ;840
            P1_P1_P2_ADS_n <= #1 1'b0; $display(";A 841");		//(= P1_P1_P2_ADS_n    0b0)) ;841
            P1_P1_P2_State <= #1 3'sb000; $display(";A 842");		//(= P1_P1_P2_State    0b000)) ;842
            P1_P1_P2_StateNA <= #1 1'b0; $display(";A 843");		//(= P1_P1_P2_StateNA    0b0)) ;843
            P1_P1_P2_StateBS16 <= #1 1'b0; $display(";A 844");		//(= P1_P1_P2_StateBS16    0b0)) ;844
            P1_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 845");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000000)) ;845
        end
        else begin
            $display(";A 835");		//(= (bv-comp P1_P1_P2_RESET  0b1)   0b0)) ;835
            case (P1_P1_P2_State)
                3'b000 :
                    begin
                        $display(";A 846");		//(= P1_P1_P2_State    0b000)) ;846
                        P1_P1_P2_D_C_n <= #1 1'b1; $display(";A 847");		//(= P1_P1_P2_D_C_n    0b1)) ;847
                        P1_P1_P2_ADS_n <= #1 1'b1; $display(";A 848");		//(= P1_P1_P2_ADS_n    0b1)) ;848
                        P1_P1_P2_State <= #1 3'sb001; $display(";A 849");		//(= P1_P1_P2_State    0b001)) ;849
                        P1_P1_P2_StateNA <= #1 1'b1; $display(";A 850");		//(= P1_P1_P2_StateNA    0b1)) ;850
                        P1_P1_P2_StateBS16 <= #1 1'b1; $display(";A 851");		//(= P1_P1_P2_StateBS16    0b1)) ;851
                        P1_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 852");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;852
                        P1_P1_P2_State <= #1 3'sb001; $display(";A 853");		//(= P1_P1_P2_State    0b001)) ;853
                    end
                3'b001 :
                    begin
                        $display(";A 854");		//(= P1_P1_P2_State    0b001)) ;854
                        if ((P1_P1_P2_RequestPending == 1'b1)) begin
                            $display(";A 855");		//(= (bv-comp P1_P1_P2_RequestPending  0b1)   0b1)) ;855
                            P1_P1_P2_State <= #1 3'sb010; $display(";A 857");		//(= P1_P1_P2_State    0b010)) ;857
                        end
                        else begin
                            $display(";A 856");		//(= (bv-comp P1_P1_P2_RequestPending  0b1)   0b0)) ;856
                            if ((P1_P1_P2_HOLD == 1'b1)) begin
                                $display(";A 858");		//(= (bv-comp P1_P1_P2_HOLD  0b1)   0b1)) ;858
                                P1_P1_P2_State <= #1 3'sb101; $display(";A 860");		//(= P1_P1_P2_State    0b101)) ;860
                            end
                            else begin
                                $display(";A 859");		//(= (bv-comp P1_P1_P2_HOLD  0b1)   0b0)) ;859
                                P1_P1_P2_State <= #1 3'sb001; $display(";A 861");		//(= P1_P1_P2_State    0b001)) ;861
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 862");		//(= P1_P1_P2_State    0b010)) ;862
                        P1_P1_P2_Address <= #1 ((P1_P1_P2_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 863");		//(= P1_P1_P2_Address    (bv-smod (bv-sdiv P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;863
                        P1_P1_P2_BE_n <= #1 P1_P1_P2_ByteEnable; $display(";A 864");		//(= P1_P1_P2_BE_n    P1_P1_P2_ByteEnable )) ;864
                        P1_P1_P2_M_IO_n <= #1 P1_P1_P2_MemoryFetch; $display(";A 865");		//(= P1_P1_P2_M_IO_n    P1_P1_P2_MemoryFetch )) ;865
                        if ((P1_P1_P2_ReadRequest == 1'b1)) begin
                            $display(";A 866");		//(= (bv-comp P1_P1_P2_ReadRequest  0b1)   0b1)) ;866
                            P1_P1_P2_W_R_n <= #1 1'b0; $display(";A 868");		//(= P1_P1_P2_W_R_n    0b0)) ;868
                        end
                        else begin
                            $display(";A 867");		//(= (bv-comp P1_P1_P2_ReadRequest  0b1)   0b0)) ;867
                            P1_P1_P2_W_R_n <= #1 1'b1; $display(";A 869");		//(= P1_P1_P2_W_R_n    0b1)) ;869
                        end
                        if ((P1_P1_P2_CodeFetch == 1'b1)) begin
                            $display(";A 870");		//(= (bv-comp P1_P1_P2_CodeFetch  0b1)   0b1)) ;870
                            P1_P1_P2_D_C_n <= #1 1'b0; $display(";A 872");		//(= P1_P1_P2_D_C_n    0b0)) ;872
                        end
                        else begin
                            $display(";A 871");		//(= (bv-comp P1_P1_P2_CodeFetch  0b1)   0b0)) ;871
                            P1_P1_P2_D_C_n <= #1 1'b1; $display(";A 873");		//(= P1_P1_P2_D_C_n    0b1)) ;873
                        end
                        P1_P1_P2_ADS_n <= #1 1'b0; $display(";A 874");		//(= P1_P1_P2_ADS_n    0b0)) ;874
                        P1_P1_P2_State <= #1 3'sb011; $display(";A 875");		//(= P1_P1_P2_State    0b011)) ;875
                    end
                3'b011 :
                    begin
                        $display(";A 876");		//(= P1_P1_P2_State    0b011)) ;876
                        if ((((P1_P1_P2_READY_n == 1'b0) & (P1_P1_P2_HOLD == 1'b0)) & (P1_P1_P2_RequestPending == 1'b1))) begin
                            $display(";A 877");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b1))   0b1)) ;877
                            P1_P1_P2_State <= #1 3'sb010; $display(";A 879");		//(= P1_P1_P2_State    0b010)) ;879
                        end
                        else begin
                            $display(";A 878");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b1))   0b0)) ;878
                            if (((P1_P1_P2_READY_n == 1'b1) & (P1_P1_P2_NA_n == 1'b1))) begin
                                $display(";A 880");		//(= (bv-and (bv-comp P1_P1_P2_READY_n  0b1) (bv-comp P1_P1_P2_NA_n  0b1))   0b1)) ;880
                            end
                            else begin
                                $display(";A 881");		//(= (bv-and (bv-comp P1_P1_P2_READY_n  0b1) (bv-comp P1_P1_P2_NA_n  0b1))   0b0)) ;881
                                if ((((P1_P1_P2_RequestPending == 1'b1) | (P1_P1_P2_HOLD == 1'b1)) & ((P1_P1_P2_READY_n == 1'b1) & (P1_P1_P2_NA_n == 1'b0)))) begin
                                    $display(";A 882");		//(= (bv-and (bv-or (bv-comp P1_P1_P2_RequestPending  0b1) (bv-comp P1_P1_P2_HOLD  0b1)) (bv-and (bv-comp P1_P1_P2_READY_n  0b1) (bv-comp P1_P1_P2_NA_n  0b0)))   0b1)) ;882
                                    P1_P1_P2_State <= #1 3'sb111; $display(";A 884");		//(= P1_P1_P2_State    0b111)) ;884
                                end
                                else begin
                                    $display(";A 883");		//(= (bv-and (bv-or (bv-comp P1_P1_P2_RequestPending  0b1) (bv-comp P1_P1_P2_HOLD  0b1)) (bv-and (bv-comp P1_P1_P2_READY_n  0b1) (bv-comp P1_P1_P2_NA_n  0b0)))   0b0)) ;883
                                    if (((((P1_P1_P2_RequestPending == 1'b1) & (P1_P1_P2_HOLD == 1'b0)) & (P1_P1_P2_READY_n == 1'b1)) & (P1_P1_P2_NA_n == 1'b0))) begin
                                        $display(";A 885");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P1_P2_RequestPending  0b1) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_READY_n  0b1)) (bv-comp P1_P1_P2_NA_n  0b0))   0b1)) ;885
                                        P1_P1_P2_State <= #1 3'sb110; $display(";A 887");		//(= P1_P1_P2_State    0b110)) ;887
                                    end
                                    else begin
                                        $display(";A 886");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P1_P2_RequestPending  0b1) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_READY_n  0b1)) (bv-comp P1_P1_P2_NA_n  0b0))   0b0)) ;886
                                        if ((((P1_P1_P2_RequestPending == 1'b0) & (P1_P1_P2_HOLD == 1'b0)) & (P1_P1_P2_READY_n == 1'b0))) begin
                                            $display(";A 888");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_RequestPending  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_READY_n  0b0))   0b1)) ;888
                                            P1_P1_P2_State <= #1 3'sb001; $display(";A 890");		//(= P1_P1_P2_State    0b001)) ;890
                                        end
                                        else begin
                                            $display(";A 889");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_RequestPending  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_READY_n  0b0))   0b0)) ;889
                                            if (((P1_P1_P2_HOLD == 1'b1) & (P1_P1_P2_READY_n == 1'b1))) begin
                                                $display(";A 891");		//(= (bv-and (bv-comp P1_P1_P2_HOLD  0b1) (bv-comp P1_P1_P2_READY_n  0b1))   0b1)) ;891
                                                P1_P1_P2_State <= #1 3'sb101; $display(";A 893");		//(= P1_P1_P2_State    0b101)) ;893
                                            end
                                            else begin
                                                $display(";A 892");		//(= (bv-and (bv-comp P1_P1_P2_HOLD  0b1) (bv-comp P1_P1_P2_READY_n  0b1))   0b0)) ;892
                                                P1_P1_P2_State <= #1 3'sb011; $display(";A 894");		//(= P1_P1_P2_State    0b011)) ;894
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P1_P1_P2_StateBS16 <= #1 P1_P1_P2_BS16_n; $display(";A 895");		//(= P1_P1_P2_StateBS16    P1_P1_P2_BS16_n )) ;895
                        if ((P1_P1_P2_BS16_n == 1'b0)) begin
                            $display(";A 896");		//(= (bv-comp P1_P1_P2_BS16_n  0b0)   0b1)) ;896
                            P1_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 898");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000001)) ;898
                        end
                        else begin
                            $display(";A 897");		//(= (bv-comp P1_P1_P2_BS16_n  0b0)   0b0)) ;897
                            P1_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 899");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;899
                        end
                        P1_P1_P2_StateNA <= #1 P1_P1_P2_NA_n; $display(";A 900");		//(= P1_P1_P2_StateNA    P1_P1_P2_NA_n )) ;900
                        P1_P1_P2_ADS_n <= #1 1'b1; $display(";A 901");		//(= P1_P1_P2_ADS_n    0b1)) ;901
                    end
                3'b100 :
                    begin
                        $display(";A 902");		//(= P1_P1_P2_State    0b100)) ;902
                        if ((((P1_P1_P2_NA_n == 1'b0) & (P1_P1_P2_HOLD == 1'b0)) & (P1_P1_P2_RequestPending == 1'b1))) begin
                            $display(";A 903");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_NA_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b1))   0b1)) ;903
                            P1_P1_P2_State <= #1 3'sb110; $display(";A 905");		//(= P1_P1_P2_State    0b110)) ;905
                        end
                        else begin
                            $display(";A 904");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_NA_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b1))   0b0)) ;904
                            if (((P1_P1_P2_NA_n == 1'b0) & ((P1_P1_P2_HOLD == 1'b1) | (P1_P1_P2_RequestPending == 1'b0)))) begin
                                $display(";A 906");		//(= (bv-and (bv-comp P1_P1_P2_NA_n  0b0) (bv-or (bv-comp P1_P1_P2_HOLD  0b1) (bv-comp P1_P1_P2_RequestPending  0b0)))   0b1)) ;906
                                P1_P1_P2_State <= #1 3'sb111; $display(";A 908");		//(= P1_P1_P2_State    0b111)) ;908
                            end
                            else begin
                                $display(";A 907");		//(= (bv-and (bv-comp P1_P1_P2_NA_n  0b0) (bv-or (bv-comp P1_P1_P2_HOLD  0b1) (bv-comp P1_P1_P2_RequestPending  0b0)))   0b0)) ;907
                                if ((P1_P1_P2_NA_n == 1'b1)) begin
                                    $display(";A 909");		//(= (bv-comp P1_P1_P2_NA_n  0b1)   0b1)) ;909
                                    P1_P1_P2_State <= #1 3'sb011; $display(";A 911");		//(= P1_P1_P2_State    0b011)) ;911
                                end
                                else begin
                                    $display(";A 910");		//(= (bv-comp P1_P1_P2_NA_n  0b1)   0b0)) ;910
                                    P1_P1_P2_State <= #1 3'sb100; $display(";A 912");		//(= P1_P1_P2_State    0b100)) ;912
                                end
                            end
                        end
                        P1_P1_P2_StateBS16 <= #1 P1_P1_P2_BS16_n; $display(";A 913");		//(= P1_P1_P2_StateBS16    P1_P1_P2_BS16_n )) ;913
                        if ((P1_P1_P2_BS16_n == 1'b0)) begin
                            $display(";A 914");		//(= (bv-comp P1_P1_P2_BS16_n  0b0)   0b1)) ;914
                            P1_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 916");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000001)) ;916
                        end
                        else begin
                            $display(";A 915");		//(= (bv-comp P1_P1_P2_BS16_n  0b0)   0b0)) ;915
                            P1_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 917");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;917
                        end
                        P1_P1_P2_StateNA <= #1 P1_P1_P2_NA_n; $display(";A 918");		//(= P1_P1_P2_StateNA    P1_P1_P2_NA_n )) ;918
                        P1_P1_P2_ADS_n <= #1 1'b1; $display(";A 919");		//(= P1_P1_P2_ADS_n    0b1)) ;919
                    end
                3'b101 :
                    begin
                        $display(";A 920");		//(= P1_P1_P2_State    0b101)) ;920
                        if (((P1_P1_P2_HOLD == 1'b0) & (P1_P1_P2_RequestPending == 1'b1))) begin
                            $display(";A 921");		//(= (bv-and (bv-comp P1_P1_P2_HOLD  0b0) (bv-comp P1_P1_P2_RequestPending  0b1))   0b1)) ;921
                            P1_P1_P2_State <= #1 3'sb010; $display(";A 923");		//(= P1_P1_P2_State    0b010)) ;923
                        end
                        else begin
                            $display(";A 922");		//(= (bv-and (bv-comp P1_P1_P2_HOLD  0b0) (bv-comp P1_P1_P2_RequestPending  0b1))   0b0)) ;922
                            if (((P1_P1_P2_HOLD == 1'b0) & (P1_P1_P2_RequestPending == 1'b0))) begin
                                $display(";A 924");		//(= (bv-and (bv-comp P1_P1_P2_HOLD  0b0) (bv-comp P1_P1_P2_RequestPending  0b0))   0b1)) ;924
                                P1_P1_P2_State <= #1 3'sb001; $display(";A 926");		//(= P1_P1_P2_State    0b001)) ;926
                            end
                            else begin
                                $display(";A 925");		//(= (bv-and (bv-comp P1_P1_P2_HOLD  0b0) (bv-comp P1_P1_P2_RequestPending  0b0))   0b0)) ;925
                                P1_P1_P2_State <= #1 3'sb101; $display(";A 927");		//(= P1_P1_P2_State    0b101)) ;927
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 928");		//(= P1_P1_P2_State    0b110)) ;928
                        P1_P1_P2_Address <= #1 ((P1_P1_P2_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 929");		//(= P1_P1_P2_Address    (bv-smod (bv-sdiv P1_P1_P2_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;929
                        P1_P1_P2_BE_n <= #1 P1_P1_P2_ByteEnable; $display(";A 930");		//(= P1_P1_P2_BE_n    P1_P1_P2_ByteEnable )) ;930
                        P1_P1_P2_M_IO_n <= #1 P1_P1_P2_MemoryFetch; $display(";A 931");		//(= P1_P1_P2_M_IO_n    P1_P1_P2_MemoryFetch )) ;931
                        if ((P1_P1_P2_ReadRequest == 1'b1)) begin
                            $display(";A 932");		//(= (bv-comp P1_P1_P2_ReadRequest  0b1)   0b1)) ;932
                            P1_P1_P2_W_R_n <= #1 1'b0; $display(";A 934");		//(= P1_P1_P2_W_R_n    0b0)) ;934
                        end
                        else begin
                            $display(";A 933");		//(= (bv-comp P1_P1_P2_ReadRequest  0b1)   0b0)) ;933
                            P1_P1_P2_W_R_n <= #1 1'b1; $display(";A 935");		//(= P1_P1_P2_W_R_n    0b1)) ;935
                        end
                        if ((P1_P1_P2_CodeFetch == 1'b1)) begin
                            $display(";A 936");		//(= (bv-comp P1_P1_P2_CodeFetch  0b1)   0b1)) ;936
                            P1_P1_P2_D_C_n <= #1 1'b0; $display(";A 938");		//(= P1_P1_P2_D_C_n    0b0)) ;938
                        end
                        else begin
                            $display(";A 937");		//(= (bv-comp P1_P1_P2_CodeFetch  0b1)   0b0)) ;937
                            P1_P1_P2_D_C_n <= #1 1'b1; $display(";A 939");		//(= P1_P1_P2_D_C_n    0b1)) ;939
                        end
                        P1_P1_P2_ADS_n <= #1 1'b0; $display(";A 940");		//(= P1_P1_P2_ADS_n    0b0)) ;940
                        if ((P1_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 941");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;941
                            P1_P1_P2_State <= #1 3'sb100; $display(";A 943");		//(= P1_P1_P2_State    0b100)) ;943
                        end
                        else begin
                            $display(";A 942");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;942
                            P1_P1_P2_State <= #1 3'sb110; $display(";A 944");		//(= P1_P1_P2_State    0b110)) ;944
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 945");		//(= P1_P1_P2_State    0b111)) ;945
                        if ((((P1_P1_P2_READY_n == 1'b1) & (P1_P1_P2_RequestPending == 1'b1)) & (P1_P1_P2_HOLD == 1'b0))) begin
                            $display(";A 946");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b1) (bv-comp P1_P1_P2_RequestPending  0b1)) (bv-comp P1_P1_P2_HOLD  0b0))   0b1)) ;946
                            P1_P1_P2_State <= #1 3'sb110; $display(";A 948");		//(= P1_P1_P2_State    0b110)) ;948
                        end
                        else begin
                            $display(";A 947");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b1) (bv-comp P1_P1_P2_RequestPending  0b1)) (bv-comp P1_P1_P2_HOLD  0b0))   0b0)) ;947
                            if (((P1_P1_P2_READY_n == 1'b0) & (P1_P1_P2_HOLD == 1'b1))) begin
                                $display(";A 949");		//(= (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b1))   0b1)) ;949
                                P1_P1_P2_State <= #1 3'sb101; $display(";A 951");		//(= P1_P1_P2_State    0b101)) ;951
                            end
                            else begin
                                $display(";A 950");		//(= (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b1))   0b0)) ;950
                                if ((((P1_P1_P2_READY_n == 1'b0) & (P1_P1_P2_HOLD == 1'b0)) & (P1_P1_P2_RequestPending == 1'b1))) begin
                                    $display(";A 952");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b1))   0b1)) ;952
                                    P1_P1_P2_State <= #1 3'sb010; $display(";A 954");		//(= P1_P1_P2_State    0b010)) ;954
                                end
                                else begin
                                    $display(";A 953");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b1))   0b0)) ;953
                                    if ((((P1_P1_P2_READY_n == 1'b0) & (P1_P1_P2_HOLD == 1'b0)) & (P1_P1_P2_RequestPending == 1'b0))) begin
                                        $display(";A 955");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b0))   0b1)) ;955
                                        P1_P1_P2_State <= #1 3'sb001; $display(";A 957");		//(= P1_P1_P2_State    0b001)) ;957
                                    end
                                    else begin
                                        $display(";A 956");		//(= (bv-and (bv-and (bv-comp P1_P1_P2_READY_n  0b0) (bv-comp P1_P1_P2_HOLD  0b0)) (bv-comp P1_P1_P2_RequestPending  0b0))   0b0)) ;956
                                        P1_P1_P2_State <= #1 3'sb111; $display(";A 958");		//(= P1_P1_P2_State    0b111)) ;958
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:1259
    always @(posedge P1_P1_P2_RESET or posedge P1_P1_P2_CLOCK) begin
        if ((P1_P1_P2_RESET == 1'b1)) begin
            $display(";A 959");		//(= (bv-comp P1_P1_P2_RESET  0b1)   0b1)) ;959
            P1_P1_P2_State2 = 4'sb0000; $display(";A 961");		//(= P1_P1_P2_State2    0b0000)) ;961
            P1_P1_P2_InstQueue[0] = 8'b00000000; $display(";A 962");		//(= P1_P1_P2_InstQueue    0b00000000)) ;962
            P1_P1_P2_InstQueue[1] = 8'b00000000; $display(";A 963");		//(= P1_P1_P2_InstQueue    0b00000000)) ;963
            P1_P1_P2_InstQueue[2] = 8'b00000000; $display(";A 964");		//(= P1_P1_P2_InstQueue    0b00000000)) ;964
            P1_P1_P2_InstQueue[3] = 8'b00000000; $display(";A 965");		//(= P1_P1_P2_InstQueue    0b00000000)) ;965
            P1_P1_P2_InstQueue[4] = 8'b00000000; $display(";A 966");		//(= P1_P1_P2_InstQueue    0b00000000)) ;966
            P1_P1_P2_InstQueue[5] = 8'b00000000; $display(";A 967");		//(= P1_P1_P2_InstQueue    0b00000000)) ;967
            P1_P1_P2_InstQueue[6] = 8'b00000000; $display(";A 968");		//(= P1_P1_P2_InstQueue    0b00000000)) ;968
            P1_P1_P2_InstQueue[7] = 8'b00000000; $display(";A 969");		//(= P1_P1_P2_InstQueue    0b00000000)) ;969
            P1_P1_P2_InstQueue[8] = 8'b00000000; $display(";A 970");		//(= P1_P1_P2_InstQueue    0b00000000)) ;970
            P1_P1_P2_InstQueue[9] = 8'b00000000; $display(";A 971");		//(= P1_P1_P2_InstQueue    0b00000000)) ;971
            P1_P1_P2_InstQueue[10] = 8'b00000000; $display(";A 972");		//(= P1_P1_P2_InstQueue    0b00000000)) ;972
            P1_P1_P2_InstQueue[11] = 8'b00000000; $display(";A 973");		//(= P1_P1_P2_InstQueue    0b00000000)) ;973
            P1_P1_P2_InstQueue[12] = 8'b00000000; $display(";A 974");		//(= P1_P1_P2_InstQueue    0b00000000)) ;974
            P1_P1_P2_InstQueue[13] = 8'b00000000; $display(";A 975");		//(= P1_P1_P2_InstQueue    0b00000000)) ;975
            P1_P1_P2_InstQueue[14] = 8'b00000000; $display(";A 976");		//(= P1_P1_P2_InstQueue    0b00000000)) ;976
            P1_P1_P2_InstQueue[15] = 8'b00000000; $display(";A 977");		//(= P1_P1_P2_InstQueue    0b00000000)) ;977
            P1_P1_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 978");		//(= P1_P1_P2_InstQueueRd_Addr    0b00000)) ;978
            P1_P1_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 979");		//(= P1_P1_P2_InstQueueWr_Addr    0b00000)) ;979
            P1_P1_P2_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 980");		//(= P1_P1_P2_InstAddrPointer    0b00000000000000000000000000000000)) ;980
            P1_P1_P2_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 981");		//(= P1_P1_P2_PhyAddrPointer    0b00000000000000000000000000000000)) ;981
            P1_P1_P2_Extended = 1'b0; $display(";A 982");		//(= P1_P1_P2_Extended    0b0)) ;982
            P1_P1_P2_More = 1'b0; $display(";A 983");		//(= P1_P1_P2_More    0b0)) ;983
            P1_P1_P2_Flush = 1'b0; $display(";A 984");		//(= P1_P1_P2_Flush    0b0)) ;984
            P1_P1_P2_lWord = 16'sb0000000000000000; $display(";A 985");		//(= P1_P1_P2_lWord    0b0000000000000000)) ;985
            P1_P1_P2_uWord = 15'sb000000000000000; $display(";A 986");		//(= P1_P1_P2_uWord    0b000000000000000)) ;986
            P1_P1_P2_fWord = 32'sb00000000000000000000000000000000; $display(";A 987");		//(= P1_P1_P2_fWord    0b00000000000000000000000000000000)) ;987
            P1_P1_P2_CodeFetch <= #1 1'b0; $display(";A 988");		//(= P1_P1_P2_CodeFetch    0b0)) ;988
            P1_P1_P2_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 989");		//(= P1_P1_P2_Datao    0b00000000000000000000000000000000)) ;989
            P1_P1_P2_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 990");		//(= P1_P1_P2_EAX    0b00000000000000000000000000000000)) ;990
            P1_P1_P2_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 991");		//(= P1_P1_P2_EBX    0b00000000000000000000000000000000)) ;991
            P1_P1_P2_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 992");		//(= P1_P1_P2_rEIP    0b00000000000000000000000000000000)) ;992
            P1_P1_P2_ReadRequest <= #1 1'b0; $display(";A 993");		//(= P1_P1_P2_ReadRequest    0b0)) ;993
            P1_P1_P2_MemoryFetch <= #1 1'b0; $display(";A 994");		//(= P1_P1_P2_MemoryFetch    0b0)) ;994
            P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 995");		//(= P1_P1_P2_RequestPending    0b0)) ;995
        end
        else begin
            $display(";A 960");		//(= (bv-comp P1_P1_P2_RESET  0b1)   0b0)) ;960
            case (P1_P1_P2_State2)
                4'b0000 :
                    begin
                        $display(";A 996");		//(= P1_P1_P2_State2    0b0000)) ;996
                        P1_P1_P2_PhyAddrPointer = P1_P1_P2_rEIP; $display(";A 997");		//(= P1_P1_P2_PhyAddrPointer    P1_P1_P2_rEIP )) ;997
                        P1_P1_P2_InstAddrPointer = P1_P1_P2_PhyAddrPointer; $display(";A 998");		//(= P1_P1_P2_InstAddrPointer    P1_P1_P2_PhyAddrPointer )) ;998
                        P1_P1_P2_State2 = 4'sb0001; $display(";A 999");		//(= P1_P1_P2_State2    0b0001)) ;999
                        P1_P1_P2_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 1000");		//(= P1_P1_P2_rEIP    0b00000000000011111111111111110000)) ;1000
                        P1_P1_P2_ReadRequest <= #1 1'b1; $display(";A 1001");		//(= P1_P1_P2_ReadRequest    0b1)) ;1001
                        P1_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 1002");		//(= P1_P1_P2_MemoryFetch    0b1)) ;1002
                        P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1003");		//(= P1_P1_P2_RequestPending    0b1)) ;1003
                    end
                4'b0001 :
                    begin
                        $display(";A 1004");		//(= P1_P1_P2_State2    0b0001)) ;1004
                        P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1005");		//(= P1_P1_P2_RequestPending    0b1)) ;1005
                        P1_P1_P2_ReadRequest <= #1 1'b1; $display(";A 1006");		//(= P1_P1_P2_ReadRequest    0b1)) ;1006
                        P1_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 1007");		//(= P1_P1_P2_MemoryFetch    0b1)) ;1007
                        P1_P1_P2_CodeFetch <= #1 1'b1; $display(";A 1008");		//(= P1_P1_P2_CodeFetch    0b1)) ;1008
                        if ((P1_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 1009");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1009
                            P1_P1_P2_State2 = 4'sb0010; $display(";A 1011");		//(= P1_P1_P2_State2    0b0010)) ;1011
                        end
                        else begin
                            $display(";A 1010");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1010
                            P1_P1_P2_State2 = 4'sb0001; $display(";A 1012");		//(= P1_P1_P2_State2    0b0001)) ;1012
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 1013");		//(= P1_P1_P2_State2    0b0010)) ;1013
                        P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1014");		//(= P1_P1_P2_RequestPending    0b0)) ;1014
                        P1_P1_P2_InstQueue[P1_P1_P2_InstQueueWr_Addr] = (P1_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 1015");		//(= P1_P1_P2_InstQueue    (bv-smod P1_P1_P2_Datai  0b00000000000000000000000100000000))) ;1015
                        P1_P1_P2_InstQueueWr_Addr = ((P1_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1016");		//(= P1_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1016
                        P1_P1_P2_InstQueue[P1_P1_P2_InstQueueWr_Addr] = (P1_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 1017");		//(= P1_P1_P2_InstQueue    (bv-smod P1_P1_P2_Datai  0b00000000000000000000000100000000))) ;1017
                        P1_P1_P2_InstQueueWr_Addr = ((P1_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1018");		//(= P1_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1018
                        if ((P1_P1_P2_StateBS16 == 1'b1)) begin
                            $display(";A 1019");		//(= (bv-comp P1_P1_P2_StateBS16  0b1)   0b1)) ;1019
                            P1_P1_P2_InstQueue[P1_P1_P2_InstQueueWr_Addr] = ((P1_P1_P2_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 1021");		//(= P1_P1_P2_InstQueue    (bv-smod (bv-sdiv P1_P1_P2_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;1021
                            P1_P1_P2_InstQueueWr_Addr = ((P1_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1022");		//(= P1_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1022
                            P1_P1_P2_InstQueue[P1_P1_P2_InstQueueWr_Addr] = ((P1_P1_P2_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 1023");		//(= P1_P1_P2_InstQueue    (bv-smod (bv-sdiv P1_P1_P2_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;1023
                            P1_P1_P2_InstQueueWr_Addr = ((P1_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1024");		//(= P1_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1024
                            P1_P1_P2_PhyAddrPointer = (P1_P1_P2_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 1025");		//(= P1_P1_P2_PhyAddrPointer    (bv-add P1_P1_P2_PhyAddrPointer  0b00000000000000000000000000000100))) ;1025
                            P1_P1_P2_State2 = 4'sb0101; $display(";A 1026");		//(= P1_P1_P2_State2    0b0101)) ;1026
                        end
                        else begin
                            $display(";A 1020");		//(= (bv-comp P1_P1_P2_StateBS16  0b1)   0b0)) ;1020
                            P1_P1_P2_PhyAddrPointer = (P1_P1_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1027");		//(= P1_P1_P2_PhyAddrPointer    (bv-add P1_P1_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;1027
                            if ((P1_P1_P2_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 1028");		//(= (bool-to-bv (bv-slt P1_P1_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;1028
                                P1_P1_P2_rEIP <= #1 (-P1_P1_P2_PhyAddrPointer); $display(";A 1030");		//(= P1_P1_P2_rEIP    (bv-neg P1_P1_P2_PhyAddrPointer ))) ;1030
                            end
                            else begin
                                $display(";A 1029");		//(= (bool-to-bv (bv-slt P1_P1_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;1029
                                P1_P1_P2_rEIP <= #1 P1_P1_P2_PhyAddrPointer; $display(";A 1031");		//(= P1_P1_P2_rEIP    P1_P1_P2_PhyAddrPointer )) ;1031
                            end
                            P1_P1_P2_State2 = 4'sb0011; $display(";A 1032");		//(= P1_P1_P2_State2    0b0011)) ;1032
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 1033");		//(= P1_P1_P2_State2    0b0011)) ;1033
                        P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1034");		//(= P1_P1_P2_RequestPending    0b1)) ;1034
                        if ((P1_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 1035");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1035
                            P1_P1_P2_State2 = 4'sb0100; $display(";A 1037");		//(= P1_P1_P2_State2    0b0100)) ;1037
                        end
                        else begin
                            $display(";A 1036");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1036
                            P1_P1_P2_State2 = 4'sb0011; $display(";A 1038");		//(= P1_P1_P2_State2    0b0011)) ;1038
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 1039");		//(= P1_P1_P2_State2    0b0100)) ;1039
                        P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1040");		//(= P1_P1_P2_RequestPending    0b0)) ;1040
                        P1_P1_P2_InstQueue[P1_P1_P2_InstQueueWr_Addr] = (P1_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 1041");		//(= P1_P1_P2_InstQueue    (bv-smod P1_P1_P2_Datai  0b00000000000000000000000100000000))) ;1041
                        P1_P1_P2_InstQueueWr_Addr = ((P1_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1042");		//(= P1_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1042
                        P1_P1_P2_InstQueue[P1_P1_P2_InstQueueWr_Addr] = (P1_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 1043");		//(= P1_P1_P2_InstQueue    (bv-smod P1_P1_P2_Datai  0b00000000000000000000000100000000))) ;1043
                        P1_P1_P2_InstQueueWr_Addr = ((P1_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1044");		//(= P1_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1044
                        P1_P1_P2_PhyAddrPointer = (P1_P1_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1045");		//(= P1_P1_P2_PhyAddrPointer    (bv-add P1_P1_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;1045
                        P1_P1_P2_State2 = 4'sb0101; $display(";A 1046");		//(= P1_P1_P2_State2    0b0101)) ;1046
                    end
                4'b0101 :
                    begin
                        $display(";A 1047");		//(= P1_P1_P2_State2    0b0101)) ;1047
                        case (P1_P1_P2_InstQueue[P1_P1_P2_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 1048");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b10010000)) ;1048
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1049");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1049
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1050");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1050
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1051");		//(= P1_P1_P2_Flush    0b0)) ;1051
                                    P1_P1_P2_More = 1'b0; $display(";A 1052");		//(= P1_P1_P2_More    0b0)) ;1052
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 1053");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b01100110)) ;1053
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1054");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1054
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1055");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1055
                                    P1_P1_P2_Extended = 1'b1; $display(";A 1056");		//(= P1_P1_P2_Extended    0b1)) ;1056
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1057");		//(= P1_P1_P2_Flush    0b0)) ;1057
                                    P1_P1_P2_More = 1'b0; $display(";A 1058");		//(= P1_P1_P2_More    0b0)) ;1058
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 1059");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b11101011)) ;1059
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 1060");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;1060
                                        if ((P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 1062");		//(= (bool-to-bv (bv-gt P1_P1_P2_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;1062
                                            P1_P1_P2_PhyAddrPointer = ((P1_P1_P2_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 1064");		//(= P1_P1_P2_PhyAddrPointer    (bv-sub (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P1_P1_P2_InstQueue 0 )))) ;1064
                                            P1_P1_P2_InstAddrPointer = P1_P1_P2_PhyAddrPointer; $display(";A 1065");		//(= P1_P1_P2_InstAddrPointer    P1_P1_P2_PhyAddrPointer )) ;1065
                                        end
                                        else begin
                                            $display(";A 1063");		//(= (bool-to-bv (bv-gt P1_P1_P2_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;1063
                                            P1_P1_P2_PhyAddrPointer = ((P1_P1_P2_InstAddrPointer + 32'b00000000000000000000000000000010) + P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 1066");		//(= P1_P1_P2_PhyAddrPointer    (bv-add (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000010) P1_P1_P2_InstQueue 0 ))) ;1066
                                            P1_P1_P2_InstAddrPointer = P1_P1_P2_PhyAddrPointer; $display(";A 1067");		//(= P1_P1_P2_InstAddrPointer    P1_P1_P2_PhyAddrPointer )) ;1067
                                        end
                                        P1_P1_P2_Flush = 1'b1; $display(";A 1068");		//(= P1_P1_P2_Flush    0b1)) ;1068
                                        P1_P1_P2_More = 1'b0; $display(";A 1069");		//(= P1_P1_P2_More    0b0)) ;1069
                                    end
                                    else begin
                                        $display(";A 1061");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;1061
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1070");		//(= P1_P1_P2_Flush    0b0)) ;1070
                                        P1_P1_P2_More = 1'b1; $display(";A 1071");		//(= P1_P1_P2_More    0b1)) ;1071
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 1072");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b11101001)) ;1072
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 1073");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;1073
                                        P1_P1_P2_PhyAddrPointer = ((P1_P1_P2_InstAddrPointer + 32'b00000000000000000000000000000101) + P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 1075");		//(= P1_P1_P2_PhyAddrPointer    (bv-add (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000101) P1_P1_P2_InstQueue 0 ))) ;1075
                                        P1_P1_P2_InstAddrPointer = P1_P1_P2_PhyAddrPointer; $display(";A 1076");		//(= P1_P1_P2_InstAddrPointer    P1_P1_P2_PhyAddrPointer )) ;1076
                                        P1_P1_P2_Flush = 1'b1; $display(";A 1077");		//(= P1_P1_P2_Flush    0b1)) ;1077
                                        P1_P1_P2_More = 1'b0; $display(";A 1078");		//(= P1_P1_P2_More    0b0)) ;1078
                                    end
                                    else begin
                                        $display(";A 1074");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;1074
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1079");		//(= P1_P1_P2_Flush    0b0)) ;1079
                                        P1_P1_P2_More = 1'b1; $display(";A 1080");		//(= P1_P1_P2_More    0b1)) ;1080
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 1081");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b11101010)) ;1081
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1082");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1082
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1083");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1083
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1084");		//(= P1_P1_P2_Flush    0b0)) ;1084
                                    P1_P1_P2_More = 1'b0; $display(";A 1085");		//(= P1_P1_P2_More    0b0)) ;1085
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 1086");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b10110000)) ;1086
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1087");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1087
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1088");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1088
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1089");		//(= P1_P1_P2_Flush    0b0)) ;1089
                                    P1_P1_P2_More = 1'b0; $display(";A 1090");		//(= P1_P1_P2_More    0b0)) ;1090
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 1091");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b10111000)) ;1091
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 1092");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;1092
                                        P1_P1_P2_EAX <= #1 ((((P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 1094");		//(= P1_P1_P2_EAX    (bv-add (bv-add (bv-add (bv-mul P1_P1_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P1_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P1_P2_InstQueue 0  0b00000000000000000000000100000000)) P1_P1_P2_InstQueue 0 ))) ;1094
                                        P1_P1_P2_More = 1'b0; $display(";A 1095");		//(= P1_P1_P2_More    0b0)) ;1095
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1096");		//(= P1_P1_P2_Flush    0b0)) ;1096
                                        P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 1097");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;1097
                                        P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 1098");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;1098
                                    end
                                    else begin
                                        $display(";A 1093");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;1093
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1099");		//(= P1_P1_P2_Flush    0b0)) ;1099
                                        P1_P1_P2_More = 1'b1; $display(";A 1100");		//(= P1_P1_P2_More    0b1)) ;1100
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 1101");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b10111011)) ;1101
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 1102");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;1102
                                        P1_P1_P2_EBX <= #1 ((((P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P1_P2_InstQueue[((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 1104");		//(= P1_P1_P2_EBX    (bv-add (bv-add (bv-add (bv-mul P1_P1_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P1_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P1_P2_InstQueue 0  0b00000000000000000000000100000000)) P1_P1_P2_InstQueue 0 ))) ;1104
                                        P1_P1_P2_More = 1'b0; $display(";A 1105");		//(= P1_P1_P2_More    0b0)) ;1105
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1106");		//(= P1_P1_P2_Flush    0b0)) ;1106
                                        P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 1107");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;1107
                                        P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 1108");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;1108
                                    end
                                    else begin
                                        $display(";A 1103");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;1103
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1109");		//(= P1_P1_P2_Flush    0b0)) ;1109
                                        P1_P1_P2_More = 1'b1; $display(";A 1110");		//(= P1_P1_P2_More    0b1)) ;1110
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 1111");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b10001011)) ;1111
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1112");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1112
                                        if ((P1_P1_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 1114");		//(= (bool-to-bv (bv-slt P1_P1_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;1114
                                            P1_P1_P2_rEIP <= #1 (-P1_P1_P2_EBX); $display(";A 1116");		//(= P1_P1_P2_rEIP    (bv-neg P1_P1_P2_EBX ))) ;1116
                                        end
                                        else begin
                                            $display(";A 1115");		//(= (bool-to-bv (bv-slt P1_P1_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;1115
                                            P1_P1_P2_rEIP <= #1 P1_P1_P2_EBX; $display(";A 1117");		//(= P1_P1_P2_rEIP    P1_P1_P2_EBX )) ;1117
                                        end
                                        P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1118");		//(= P1_P1_P2_RequestPending    0b1)) ;1118
                                        P1_P1_P2_ReadRequest <= #1 1'b1; $display(";A 1119");		//(= P1_P1_P2_ReadRequest    0b1)) ;1119
                                        P1_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 1120");		//(= P1_P1_P2_MemoryFetch    0b1)) ;1120
                                        P1_P1_P2_CodeFetch <= #1 1'b0; $display(";A 1121");		//(= P1_P1_P2_CodeFetch    0b0)) ;1121
                                        if ((P1_P1_P2_READY_n == 1'b0)) begin
                                            $display(";A 1122");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1122
                                            P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1124");		//(= P1_P1_P2_RequestPending    0b0)) ;1124
                                            P1_P1_P2_uWord = (P1_P1_P2_Datai % 32'b00000000000000001000000000000000); $display(";A 1125");		//(= P1_P1_P2_uWord    (bv-smod P1_P1_P2_Datai  0b00000000000000001000000000000000))) ;1125
                                            if ((P1_P1_P2_StateBS16 == 1'b1)) begin
                                                $display(";A 1126");		//(= (bv-comp P1_P1_P2_StateBS16  0b1)   0b1)) ;1126
                                                P1_P1_P2_lWord = (P1_P1_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 1128");		//(= P1_P1_P2_lWord    (bv-smod P1_P1_P2_Datai  0b00000000000000010000000000000000))) ;1128
                                            end
                                            else begin
                                                $display(";A 1127");		//(= (bv-comp P1_P1_P2_StateBS16  0b1)   0b0)) ;1127
                                                P1_P1_P2_rEIP <= #1 (P1_P1_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 1129");		//(= P1_P1_P2_rEIP    (bv-add P1_P1_P2_rEIP  0b00000000000000000000000000000010))) ;1129
                                                P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1130");		//(= P1_P1_P2_RequestPending    0b1)) ;1130
                                                if ((P1_P1_P2_READY_n == 1'b0)) begin
                                                    $display(";A 1131");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1131
                                                    P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1133");		//(= P1_P1_P2_RequestPending    0b0)) ;1133
                                                    P1_P1_P2_lWord = (P1_P1_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 1134");		//(= P1_P1_P2_lWord    (bv-smod P1_P1_P2_Datai  0b00000000000000010000000000000000))) ;1134
                                                end
                                                else begin
                                                    $display(";A 1132");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1132
                                                end
                                            end
                                            if ((P1_P1_P2_READY_n == 1'b0)) begin
                                                $display(";A 1135");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1135
                                                P1_P1_P2_EAX <= #1 ((P1_P1_P2_uWord * 32'b00000000000000010000000000000000) + P1_P1_P2_lWord); $display(";A 1137");		//(= P1_P1_P2_EAX    (bv-add (bv-mul P1_P1_P2_uWord  0b00000000000000010000000000000000) P1_P1_P2_lWord ))) ;1137
                                                P1_P1_P2_More = 1'b0; $display(";A 1138");		//(= P1_P1_P2_More    0b0)) ;1138
                                                P1_P1_P2_Flush = 1'b0; $display(";A 1139");		//(= P1_P1_P2_Flush    0b0)) ;1139
                                                P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1140");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;1140
                                                P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1141");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1141
                                            end
                                            else begin
                                                $display(";A 1136");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1136
                                            end
                                        end
                                        else begin
                                            $display(";A 1123");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1123
                                        end
                                    end
                                    else begin
                                        $display(";A 1113");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1113
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1142");		//(= P1_P1_P2_Flush    0b0)) ;1142
                                        P1_P1_P2_More = 1'b1; $display(";A 1143");		//(= P1_P1_P2_More    0b1)) ;1143
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 1144");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b10001001)) ;1144
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1145");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1145
                                        if ((P1_P1_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 1147");		//(= (bool-to-bv (bv-slt P1_P1_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;1147
                                            P1_P1_P2_rEIP <= #1 P1_P1_P2_EBX; $display(";A 1149");		//(= P1_P1_P2_rEIP    P1_P1_P2_EBX )) ;1149
                                        end
                                        else begin
                                            $display(";A 1148");		//(= (bool-to-bv (bv-slt P1_P1_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;1148
                                            P1_P1_P2_rEIP <= #1 P1_P1_P2_EBX; $display(";A 1150");		//(= P1_P1_P2_rEIP    P1_P1_P2_EBX )) ;1150
                                        end
                                        P1_P1_P2_lWord = (P1_P1_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 1151");		//(= P1_P1_P2_lWord    (bv-smod P1_P1_P2_EAX  0b00000000000000010000000000000000))) ;1151
                                        P1_P1_P2_uWord = ((P1_P1_P2_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 1152");		//(= P1_P1_P2_uWord    (bv-smod (bv-sdiv P1_P1_P2_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;1152
                                        P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1153");		//(= P1_P1_P2_RequestPending    0b1)) ;1153
                                        P1_P1_P2_ReadRequest <= #1 1'b0; $display(";A 1154");		//(= P1_P1_P2_ReadRequest    0b0)) ;1154
                                        P1_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 1155");		//(= P1_P1_P2_MemoryFetch    0b1)) ;1155
                                        P1_P1_P2_CodeFetch <= #1 1'b0; $display(";A 1156");		//(= P1_P1_P2_CodeFetch    0b0)) ;1156
                                        if (((P1_P1_P2_State == 32'b00000000000000000000000000000010) | (P1_P1_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 1157");		//(= (bv-or (bv-comp P1_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P2_State  0b00000000000000000000000000000100))   0b1)) ;1157
                                            P1_P1_P2_Datao <= #1 ((P1_P1_P2_uWord * 32'b00000000000000010000000000000000) + P1_P1_P2_lWord); $display(";A 1159");		//(= P1_P1_P2_Datao    (bv-add (bv-mul P1_P1_P2_uWord  0b00000000000000010000000000000000) P1_P1_P2_lWord ))) ;1159
                                            if ((P1_P1_P2_READY_n == 1'b0)) begin
                                                $display(";A 1160");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1160
                                                P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1162");		//(= P1_P1_P2_RequestPending    0b0)) ;1162
                                                if ((P1_P1_P2_StateBS16 == 1'b0)) begin
                                                    $display(";A 1163");		//(= (bv-comp P1_P1_P2_StateBS16  0b0)   0b1)) ;1163
                                                    P1_P1_P2_rEIP <= #1 (P1_P1_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 1165");		//(= P1_P1_P2_rEIP    (bv-add P1_P1_P2_rEIP  0b00000000000000000000000000000010))) ;1165
                                                    P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1166");		//(= P1_P1_P2_RequestPending    0b1)) ;1166
                                                    P1_P1_P2_ReadRequest <= #1 1'b0; $display(";A 1167");		//(= P1_P1_P2_ReadRequest    0b0)) ;1167
                                                    P1_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 1168");		//(= P1_P1_P2_MemoryFetch    0b1)) ;1168
                                                    P1_P1_P2_CodeFetch <= #1 1'b0; $display(";A 1169");		//(= P1_P1_P2_CodeFetch    0b0)) ;1169
                                                    P1_P1_P2_State2 = 4'sb0110; $display(";A 1170");		//(= P1_P1_P2_State2    0b0110)) ;1170
                                                end
                                                else begin
                                                    $display(";A 1164");		//(= (bv-comp P1_P1_P2_StateBS16  0b0)   0b0)) ;1164
                                                end
                                                P1_P1_P2_More = 1'b0; $display(";A 1171");		//(= P1_P1_P2_More    0b0)) ;1171
                                                P1_P1_P2_Flush = 1'b0; $display(";A 1172");		//(= P1_P1_P2_Flush    0b0)) ;1172
                                                P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1173");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;1173
                                                P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1174");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1174
                                            end
                                            else begin
                                                $display(";A 1161");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1161
                                            end
                                        end
                                        else begin
                                            $display(";A 1158");		//(= (bv-or (bv-comp P1_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P2_State  0b00000000000000000000000000000100))   0b0)) ;1158
                                        end
                                    end
                                    else begin
                                        $display(";A 1146");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1146
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1175");		//(= P1_P1_P2_Flush    0b0)) ;1175
                                        P1_P1_P2_More = 1'b1; $display(";A 1176");		//(= P1_P1_P2_More    0b1)) ;1176
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 1177");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b11100100)) ;1177
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1178");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1178
                                        P1_P1_P2_rEIP <= #1 (P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 1180");		//(= P1_P1_P2_rEIP    (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;1180
                                        P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1181");		//(= P1_P1_P2_RequestPending    0b1)) ;1181
                                        P1_P1_P2_ReadRequest <= #1 1'b1; $display(";A 1182");		//(= P1_P1_P2_ReadRequest    0b1)) ;1182
                                        P1_P1_P2_MemoryFetch <= #1 1'b0; $display(";A 1183");		//(= P1_P1_P2_MemoryFetch    0b0)) ;1183
                                        P1_P1_P2_CodeFetch <= #1 1'b0; $display(";A 1184");		//(= P1_P1_P2_CodeFetch    0b0)) ;1184
                                        if ((P1_P1_P2_READY_n == 1'b0)) begin
                                            $display(";A 1185");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1185
                                            P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1187");		//(= P1_P1_P2_RequestPending    0b0)) ;1187
                                            P1_P1_P2_EAX <= #1 P1_P1_P2_Datai; $display(";A 1188");		//(= P1_P1_P2_EAX    P1_P1_P2_Datai )) ;1188
                                            P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1189");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;1189
                                            P1_P1_P2_InstQueueRd_Addr = (P1_P1_P2_InstQueueRd_Addr + 5'b00010); $display(";A 1190");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-add P1_P1_P2_InstQueueRd_Addr  0b00010))) ;1190
                                            P1_P1_P2_Flush = 1'b0; $display(";A 1191");		//(= P1_P1_P2_Flush    0b0)) ;1191
                                            P1_P1_P2_More = 1'b0; $display(";A 1192");		//(= P1_P1_P2_More    0b0)) ;1192
                                        end
                                        else begin
                                            $display(";A 1186");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1186
                                        end
                                    end
                                    else begin
                                        $display(";A 1179");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1179
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1193");		//(= P1_P1_P2_Flush    0b0)) ;1193
                                        P1_P1_P2_More = 1'b1; $display(";A 1194");		//(= P1_P1_P2_More    0b1)) ;1194
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 1195");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b11100110)) ;1195
                                    if (((P1_P1_P2_InstQueueWr_Addr - P1_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1196");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1196
                                        P1_P1_P2_rEIP <= #1 (P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 1198");		//(= P1_P1_P2_rEIP    (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;1198
                                        P1_P1_P2_RequestPending <= #1 1'b1; $display(";A 1199");		//(= P1_P1_P2_RequestPending    0b1)) ;1199
                                        P1_P1_P2_ReadRequest <= #1 1'b0; $display(";A 1200");		//(= P1_P1_P2_ReadRequest    0b0)) ;1200
                                        P1_P1_P2_MemoryFetch <= #1 1'b0; $display(";A 1201");		//(= P1_P1_P2_MemoryFetch    0b0)) ;1201
                                        P1_P1_P2_CodeFetch <= #1 1'b0; $display(";A 1202");		//(= P1_P1_P2_CodeFetch    0b0)) ;1202
                                        if (((P1_P1_P2_State == 32'b00000000000000000000000000000010) | (P1_P1_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 1203");		//(= (bv-or (bv-comp P1_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P2_State  0b00000000000000000000000000000100))   0b1)) ;1203
                                            P1_P1_P2_fWord = (P1_P1_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 1205");		//(= P1_P1_P2_fWord    (bv-smod P1_P1_P2_EAX  0b00000000000000010000000000000000))) ;1205
                                            P1_P1_P2_Datao <= #1 P1_P1_P2_fWord; $display(";A 1206");		//(= P1_P1_P2_Datao    P1_P1_P2_fWord )) ;1206
                                            if ((P1_P1_P2_READY_n == 1'b0)) begin
                                                $display(";A 1207");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1207
                                                P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1209");		//(= P1_P1_P2_RequestPending    0b0)) ;1209
                                                P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1210");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;1210
                                                P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1211");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1211
                                                P1_P1_P2_Flush = 1'b0; $display(";A 1212");		//(= P1_P1_P2_Flush    0b0)) ;1212
                                                P1_P1_P2_More = 1'b0; $display(";A 1213");		//(= P1_P1_P2_More    0b0)) ;1213
                                            end
                                            else begin
                                                $display(";A 1208");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1208
                                            end
                                        end
                                        else begin
                                            $display(";A 1204");		//(= (bv-or (bv-comp P1_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P2_State  0b00000000000000000000000000000100))   0b0)) ;1204
                                        end
                                    end
                                    else begin
                                        $display(";A 1197");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P2_InstQueueWr_Addr  P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1197
                                        P1_P1_P2_Flush = 1'b0; $display(";A 1214");		//(= P1_P1_P2_Flush    0b0)) ;1214
                                        P1_P1_P2_More = 1'b1; $display(";A 1215");		//(= P1_P1_P2_More    0b1)) ;1215
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 1216");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b00000100)) ;1216
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1217");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1217
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1218");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1218
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1219");		//(= P1_P1_P2_Flush    0b0)) ;1219
                                    P1_P1_P2_More = 1'b0; $display(";A 1220");		//(= P1_P1_P2_More    0b0)) ;1220
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 1221");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b00000101)) ;1221
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1222");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1222
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1223");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1223
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1224");		//(= P1_P1_P2_Flush    0b0)) ;1224
                                    P1_P1_P2_More = 1'b0; $display(";A 1225");		//(= P1_P1_P2_More    0b0)) ;1225
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 1226");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b11010000)) ;1226
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1227");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;1227
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1228");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1228
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1229");		//(= P1_P1_P2_Flush    0b0)) ;1229
                                    P1_P1_P2_More = 1'b0; $display(";A 1230");		//(= P1_P1_P2_More    0b0)) ;1230
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 1231");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b11000000)) ;1231
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1232");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;1232
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1233");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1233
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1234");		//(= P1_P1_P2_Flush    0b0)) ;1234
                                    P1_P1_P2_More = 1'b0; $display(";A 1235");		//(= P1_P1_P2_More    0b0)) ;1235
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 1236");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b01000000)) ;1236
                                    P1_P1_P2_EAX <= #1 (P1_P1_P2_EAX + 32'sb00000000000000000000000000000001); $display(";A 1237");		//(= P1_P1_P2_EAX    (bv-add P1_P1_P2_EAX  0b00000000000000000000000000000001))) ;1237
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1238");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1238
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1239");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1239
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1240");		//(= P1_P1_P2_Flush    0b0)) ;1240
                                    P1_P1_P2_More = 1'b0; $display(";A 1241");		//(= P1_P1_P2_More    0b0)) ;1241
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 1242");		//(= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr )   0b01000011)) ;1242
                                    P1_P1_P2_EBX <= #1 (P1_P1_P2_EBX + 32'sb00000000000000000000000000000001); $display(";A 1243");		//(= P1_P1_P2_EBX    (bv-add P1_P1_P2_EBX  0b00000000000000000000000000000001))) ;1243
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1244");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1244
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1245");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1245
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1246");		//(= P1_P1_P2_Flush    0b0)) ;1246
                                    P1_P1_P2_More = 1'b0; $display(";A 1247");		//(= P1_P1_P2_More    0b0)) ;1247
                                end
                            default:
                                begin
                                    $display(";A 1248");		//(= (and (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b10010000) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b01100110) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b11101011) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b11101001) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b11101010) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b10110000) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b10111000) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b10111011) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b10001011) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b10001001) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b11100100) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b11100110) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b00000100) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b00000101) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b11010000) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b11000000) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b01000000) (/= ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ) 0b01000011))   true)) ;1248
                                    P1_P1_P2_InstAddrPointer = (P1_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1249");		//(= P1_P1_P2_InstAddrPointer    (bv-add P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;1249
                                    P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1250");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1250
                                    P1_P1_P2_Flush = 1'b0; $display(";A 1251");		//(= P1_P1_P2_Flush    0b0)) ;1251
                                    P1_P1_P2_More = 1'b0; $display(";A 1252");		//(= P1_P1_P2_More    0b0)) ;1252
                                end
                        endcase
                        if (((~(P1_P1_P2_InstQueueRd_Addr < P1_P1_P2_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P1_P1_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P1_P1_P2_Flush) | P1_P1_P2_More))) begin
                            $display(";A 1253");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P1_P2_InstQueueRd_Addr  P1_P1_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P1_P2_Flush ) P1_P1_P2_More ))   0b1)) ;1253
                            P1_P1_P2_State2 = 4'sb0111; $display(";A 1255");		//(= P1_P1_P2_State2    0b0111)) ;1255
                        end
                        else begin
                            $display(";A 1254");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P1_P2_InstQueueRd_Addr  P1_P1_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P1_P2_Flush ) P1_P1_P2_More ))   0b0)) ;1254
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 1256");		//(= P1_P1_P2_State2    0b0110)) ;1256
                        P1_P1_P2_Datao <= #1 ((P1_P1_P2_uWord * 32'b00000000000000010000000000000000) + P1_P1_P2_lWord); $display(";A 1257");		//(= P1_P1_P2_Datao    (bv-add (bv-mul P1_P1_P2_uWord  0b00000000000000010000000000000000) P1_P1_P2_lWord ))) ;1257
                        if ((P1_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 1258");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b1)) ;1258
                            P1_P1_P2_RequestPending <= #1 1'b0; $display(";A 1260");		//(= P1_P1_P2_RequestPending    0b0)) ;1260
                            P1_P1_P2_State2 = 4'sb0101; $display(";A 1261");		//(= P1_P1_P2_State2    0b0101)) ;1261
                        end
                        else begin
                            $display(";A 1259");		//(= (bv-comp P1_P1_P2_READY_n  0b0)   0b0)) ;1259
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 1262");		//(= P1_P1_P2_State2    0b0111)) ;1262
                        if (P1_P1_P2_Flush) begin
                            $display(";A 1263");		//(= P1_P1_P2_Flush    0b1)) ;1263
                            P1_P1_P2_InstQueueRd_Addr = 5'sb00001; $display(";A 1265");		//(= P1_P1_P2_InstQueueRd_Addr    0b00001)) ;1265
                            P1_P1_P2_InstQueueWr_Addr = 5'sb00001; $display(";A 1266");		//(= P1_P1_P2_InstQueueWr_Addr    0b00001)) ;1266
                            if ((P1_P1_P2_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 1267");		//(= (bool-to-bv (bv-slt P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;1267
                                P1_P1_P2_fWord = (-P1_P1_P2_InstAddrPointer); $display(";A 1269");		//(= P1_P1_P2_fWord    (bv-neg P1_P1_P2_InstAddrPointer ))) ;1269
                            end
                            else begin
                                $display(";A 1268");		//(= (bool-to-bv (bv-slt P1_P1_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;1268
                                P1_P1_P2_fWord = P1_P1_P2_InstAddrPointer; $display(";A 1270");		//(= P1_P1_P2_fWord    P1_P1_P2_InstAddrPointer )) ;1270
                            end
                            if (((P1_P1_P2_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 1271");		//(= (bv-comp (bv-smod P1_P1_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;1271
                                P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + (P1_P1_P2_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 1273");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  (bv-smod P1_P1_P2_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;1273
                            end
                            else begin
                                $display(";A 1272");		//(= (bv-comp (bv-smod P1_P1_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;1272
                            end
                        end
                        else begin
                            $display(";A 1264");		//(= P1_P1_P2_Flush    0b0)) ;1264
                        end
                        if (((32'b00000000000000000000000000001111 - P1_P1_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 1274");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;1274
                            P1_P1_P2_State2 = 4'sb1000; $display(";A 1276");		//(= P1_P1_P2_State2    0b1000)) ;1276
                            P1_P1_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 1277");		//(= P1_P1_P2_InstQueueWr_Addr    0b00000)) ;1277
                        end
                        else begin
                            $display(";A 1275");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;1275
                            P1_P1_P2_State2 = 4'sb1001; $display(";A 1278");		//(= P1_P1_P2_State2    0b1001)) ;1278
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 1279");		//(= P1_P1_P2_State2    0b1000)) ;1279
                        if ((P1_P1_P2_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 1280");		//(= (bool-to-bv (bv-le P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;1280
                            P1_P1_P2_InstQueue[P1_P1_P2_InstQueueWr_Addr] = P1_P1_P2_InstQueue[P1_P1_P2_InstQueueRd_Addr]; $display(";A 1282");		//(= P1_P1_P2_InstQueue    ( P1_P1_P2_InstQueue P1_P1_P2_InstQueueRd_Addr ))) ;1282
                            P1_P1_P2_InstQueueRd_Addr = ((P1_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1283");		//(= P1_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1283
                            P1_P1_P2_InstQueueWr_Addr = ((P1_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1284");		//(= P1_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1284
                            P1_P1_P2_State2 = 4'sb1000; $display(";A 1285");		//(= P1_P1_P2_State2    0b1000)) ;1285
                        end
                        else begin
                            $display(";A 1281");		//(= (bool-to-bv (bv-le P1_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;1281
                            P1_P1_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 1286");		//(= P1_P1_P2_InstQueueRd_Addr    0b00000)) ;1286
                            P1_P1_P2_State2 = 4'sb1001; $display(";A 1287");		//(= P1_P1_P2_State2    0b1001)) ;1287
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 1288");		//(= P1_P1_P2_State2    0b1001)) ;1288
                        P1_P1_P2_rEIP <= #1 P1_P1_P2_PhyAddrPointer; $display(";A 1289");		//(= P1_P1_P2_rEIP    P1_P1_P2_PhyAddrPointer )) ;1289
                        P1_P1_P2_State2 = 4'sb0001; $display(";A 1290");		//(= P1_P1_P2_State2    0b0001)) ;1290
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:1698
    always @(posedge P1_P1_P2_RESET or posedge P1_P1_P2_CLOCK) begin
        if ((P1_P1_P2_RESET == 1'b1)) begin
            $display(";A 1291");		//(= (bv-comp P1_P1_P2_RESET  0b1)   0b1)) ;1291
            P1_P1_P2_ByteEnable <= #1 4'b0000; $display(";A 1293");		//(= P1_P1_P2_ByteEnable    0b0000)) ;1293
            P1_P1_P2_NonAligned <= #1 1'b0; $display(";A 1294");		//(= P1_P1_P2_NonAligned    0b0)) ;1294
        end
        else begin
            $display(";A 1292");		//(= (bv-comp P1_P1_P2_RESET  0b1)   0b0)) ;1292
            case (P1_P1_P2_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 1295");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000000)) ;1295
                        case ((P1_P1_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 1296");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;1296
                                    P1_P1_P2_ByteEnable <= #1 4'b1110; $display(";A 1297");		//(= P1_P1_P2_ByteEnable    0b1110)) ;1297
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 1298");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;1298
                                    P1_P1_P2_ByteEnable <= #1 4'b1101; $display(";A 1299");		//(= P1_P1_P2_ByteEnable    0b1101)) ;1299
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 1300");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;1300
                                    P1_P1_P2_ByteEnable <= #1 4'b1011; $display(";A 1301");		//(= P1_P1_P2_ByteEnable    0b1011)) ;1301
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 1302");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;1302
                                    P1_P1_P2_ByteEnable <= #1 4'b0111; $display(";A 1303");		//(= P1_P1_P2_ByteEnable    0b0111)) ;1303
                                end
                            default:
                                begin
                                    $display(";A 1304");		//(= (and (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;1304
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 1305");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000001)) ;1305
                        case ((P1_P1_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 1306");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;1306
                                    P1_P1_P2_ByteEnable <= #1 4'b1100; $display(";A 1307");		//(= P1_P1_P2_ByteEnable    0b1100)) ;1307
                                    P1_P1_P2_NonAligned <= #1 1'b0; $display(";A 1308");		//(= P1_P1_P2_NonAligned    0b0)) ;1308
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 1309");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;1309
                                    P1_P1_P2_ByteEnable <= #1 4'b1001; $display(";A 1310");		//(= P1_P1_P2_ByteEnable    0b1001)) ;1310
                                    P1_P1_P2_NonAligned <= #1 1'b0; $display(";A 1311");		//(= P1_P1_P2_NonAligned    0b0)) ;1311
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 1312");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;1312
                                    P1_P1_P2_ByteEnable <= #1 4'b0011; $display(";A 1313");		//(= P1_P1_P2_ByteEnable    0b0011)) ;1313
                                    P1_P1_P2_NonAligned <= #1 1'b0; $display(";A 1314");		//(= P1_P1_P2_NonAligned    0b0)) ;1314
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 1315");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;1315
                                    P1_P1_P2_ByteEnable <= #1 4'b0111; $display(";A 1316");		//(= P1_P1_P2_ByteEnable    0b0111)) ;1316
                                    P1_P1_P2_NonAligned <= #1 1'b1; $display(";A 1317");		//(= P1_P1_P2_NonAligned    0b1)) ;1317
                                end
                            default:
                                begin
                                    $display(";A 1318");		//(= (and (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;1318
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 1319");		//(= P1_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;1319
                        case ((P1_P1_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 1320");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;1320
                                    P1_P1_P2_ByteEnable <= #1 4'b0000; $display(";A 1321");		//(= P1_P1_P2_ByteEnable    0b0000)) ;1321
                                    P1_P1_P2_NonAligned <= #1 1'b0; $display(";A 1322");		//(= P1_P1_P2_NonAligned    0b0)) ;1322
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 1323");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;1323
                                    P1_P1_P2_ByteEnable <= #1 4'b0001; $display(";A 1324");		//(= P1_P1_P2_ByteEnable    0b0001)) ;1324
                                    P1_P1_P2_NonAligned <= #1 1'b1; $display(";A 1325");		//(= P1_P1_P2_NonAligned    0b1)) ;1325
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 1326");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;1326
                                    P1_P1_P2_NonAligned <= #1 1'b1; $display(";A 1327");		//(= P1_P1_P2_NonAligned    0b1)) ;1327
                                    P1_P1_P2_ByteEnable <= #1 4'b0011; $display(";A 1328");		//(= P1_P1_P2_ByteEnable    0b0011)) ;1328
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 1329");		//(= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;1329
                                    P1_P1_P2_NonAligned <= #1 1'b1; $display(";A 1330");		//(= P1_P1_P2_NonAligned    0b1)) ;1330
                                    P1_P1_P2_ByteEnable <= #1 4'b0111; $display(";A 1331");		//(= P1_P1_P2_ByteEnable    0b0111)) ;1331
                                end
                            default:
                                begin
                                    $display(";A 1332");		//(= (and (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;1332
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 1333");		//(= (and (/= P1_P1_P2_DataWidth  0b00000000000000000000000000000000) (/= P1_P1_P2_DataWidth  0b00000000000000000000000000000001) (/= P1_P1_P2_DataWidth  0b00000000000000000000000000000010))   true)) ;1333
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:1886
    always @(posedge P1_P1_P3_RESET or posedge P1_P1_P3_CLOCK) begin
        if ((P1_P1_P3_RESET == 1'b1)) begin
            $display(";A 1334");		//(= (bv-comp P1_P1_P3_RESET  0b1)   0b1)) ;1334
            P1_P1_P3_BE_n <= #1 4'b0000; $display(";A 1336");		//(= P1_P1_P3_BE_n    0b0000)) ;1336
            P1_P1_P3_Address <= #1 30'sb000000000000000000000000000000; $display(";A 1337");		//(= P1_P1_P3_Address    0b000000000000000000000000000000)) ;1337
            P1_P1_P3_W_R_n <= #1 1'b0; $display(";A 1338");		//(= P1_P1_P3_W_R_n    0b0)) ;1338
            P1_P1_P3_D_C_n <= #1 1'b0; $display(";A 1339");		//(= P1_P1_P3_D_C_n    0b0)) ;1339
            P1_P1_P3_M_IO_n <= #1 1'b0; $display(";A 1340");		//(= P1_P1_P3_M_IO_n    0b0)) ;1340
            P1_P1_P3_ADS_n <= #1 1'b0; $display(";A 1341");		//(= P1_P1_P3_ADS_n    0b0)) ;1341
            P1_P1_P3_State <= #1 3'sb000; $display(";A 1342");		//(= P1_P1_P3_State    0b000)) ;1342
            P1_P1_P3_StateNA <= #1 1'b0; $display(";A 1343");		//(= P1_P1_P3_StateNA    0b0)) ;1343
            P1_P1_P3_StateBS16 <= #1 1'b0; $display(";A 1344");		//(= P1_P1_P3_StateBS16    0b0)) ;1344
            P1_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 1345");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000000)) ;1345
        end
        else begin
            $display(";A 1335");		//(= (bv-comp P1_P1_P3_RESET  0b1)   0b0)) ;1335
            case (P1_P1_P3_State)
                3'b000 :
                    begin
                        $display(";A 1346");		//(= P1_P1_P3_State    0b000)) ;1346
                        P1_P1_P3_D_C_n <= #1 1'b1; $display(";A 1347");		//(= P1_P1_P3_D_C_n    0b1)) ;1347
                        P1_P1_P3_ADS_n <= #1 1'b1; $display(";A 1348");		//(= P1_P1_P3_ADS_n    0b1)) ;1348
                        P1_P1_P3_State <= #1 3'sb001; $display(";A 1349");		//(= P1_P1_P3_State    0b001)) ;1349
                        P1_P1_P3_StateNA <= #1 1'b1; $display(";A 1350");		//(= P1_P1_P3_StateNA    0b1)) ;1350
                        P1_P1_P3_StateBS16 <= #1 1'b1; $display(";A 1351");		//(= P1_P1_P3_StateBS16    0b1)) ;1351
                        P1_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 1352");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;1352
                        P1_P1_P3_State <= #1 3'sb001; $display(";A 1353");		//(= P1_P1_P3_State    0b001)) ;1353
                    end
                3'b001 :
                    begin
                        $display(";A 1354");		//(= P1_P1_P3_State    0b001)) ;1354
                        if ((P1_P1_P3_RequestPending == 1'b1)) begin
                            $display(";A 1355");		//(= (bv-comp P1_P1_P3_RequestPending  0b1)   0b1)) ;1355
                            P1_P1_P3_State <= #1 3'sb010; $display(";A 1357");		//(= P1_P1_P3_State    0b010)) ;1357
                        end
                        else begin
                            $display(";A 1356");		//(= (bv-comp P1_P1_P3_RequestPending  0b1)   0b0)) ;1356
                            if ((P1_P1_P3_HOLD == 1'b1)) begin
                                $display(";A 1358");		//(= (bv-comp P1_P1_P3_HOLD  0b1)   0b1)) ;1358
                                P1_P1_P3_State <= #1 3'sb101; $display(";A 1360");		//(= P1_P1_P3_State    0b101)) ;1360
                            end
                            else begin
                                $display(";A 1359");		//(= (bv-comp P1_P1_P3_HOLD  0b1)   0b0)) ;1359
                                P1_P1_P3_State <= #1 3'sb001; $display(";A 1361");		//(= P1_P1_P3_State    0b001)) ;1361
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 1362");		//(= P1_P1_P3_State    0b010)) ;1362
                        P1_P1_P3_Address <= #1 ((P1_P1_P3_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 1363");		//(= P1_P1_P3_Address    (bv-smod (bv-sdiv P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;1363
                        P1_P1_P3_BE_n <= #1 P1_P1_P3_ByteEnable; $display(";A 1364");		//(= P1_P1_P3_BE_n    P1_P1_P3_ByteEnable )) ;1364
                        P1_P1_P3_M_IO_n <= #1 P1_P1_P3_MemoryFetch; $display(";A 1365");		//(= P1_P1_P3_M_IO_n    P1_P1_P3_MemoryFetch )) ;1365
                        if ((P1_P1_P3_ReadRequest == 1'b1)) begin
                            $display(";A 1366");		//(= (bv-comp P1_P1_P3_ReadRequest  0b1)   0b1)) ;1366
                            P1_P1_P3_W_R_n <= #1 1'b0; $display(";A 1368");		//(= P1_P1_P3_W_R_n    0b0)) ;1368
                        end
                        else begin
                            $display(";A 1367");		//(= (bv-comp P1_P1_P3_ReadRequest  0b1)   0b0)) ;1367
                            P1_P1_P3_W_R_n <= #1 1'b1; $display(";A 1369");		//(= P1_P1_P3_W_R_n    0b1)) ;1369
                        end
                        if ((P1_P1_P3_CodeFetch == 1'b1)) begin
                            $display(";A 1370");		//(= (bv-comp P1_P1_P3_CodeFetch  0b1)   0b1)) ;1370
                            P1_P1_P3_D_C_n <= #1 1'b0; $display(";A 1372");		//(= P1_P1_P3_D_C_n    0b0)) ;1372
                        end
                        else begin
                            $display(";A 1371");		//(= (bv-comp P1_P1_P3_CodeFetch  0b1)   0b0)) ;1371
                            P1_P1_P3_D_C_n <= #1 1'b1; $display(";A 1373");		//(= P1_P1_P3_D_C_n    0b1)) ;1373
                        end
                        P1_P1_P3_ADS_n <= #1 1'b0; $display(";A 1374");		//(= P1_P1_P3_ADS_n    0b0)) ;1374
                        P1_P1_P3_State <= #1 3'sb011; $display(";A 1375");		//(= P1_P1_P3_State    0b011)) ;1375
                    end
                3'b011 :
                    begin
                        $display(";A 1376");		//(= P1_P1_P3_State    0b011)) ;1376
                        if ((((P1_P1_P3_READY_n == 1'b0) & (P1_P1_P3_HOLD == 1'b0)) & (P1_P1_P3_RequestPending == 1'b1))) begin
                            $display(";A 1377");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b1))   0b1)) ;1377
                            P1_P1_P3_State <= #1 3'sb010; $display(";A 1379");		//(= P1_P1_P3_State    0b010)) ;1379
                        end
                        else begin
                            $display(";A 1378");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b1))   0b0)) ;1378
                            if (((P1_P1_P3_READY_n == 1'b1) & (P1_P1_P3_NA_n == 1'b1))) begin
                                $display(";A 1380");		//(= (bv-and (bv-comp P1_P1_P3_READY_n  0b1) (bv-comp P1_P1_P3_NA_n  0b1))   0b1)) ;1380
                            end
                            else begin
                                $display(";A 1381");		//(= (bv-and (bv-comp P1_P1_P3_READY_n  0b1) (bv-comp P1_P1_P3_NA_n  0b1))   0b0)) ;1381
                                if ((((P1_P1_P3_RequestPending == 1'b1) | (P1_P1_P3_HOLD == 1'b1)) & ((P1_P1_P3_READY_n == 1'b1) & (P1_P1_P3_NA_n == 1'b0)))) begin
                                    $display(";A 1382");		//(= (bv-and (bv-or (bv-comp P1_P1_P3_RequestPending  0b1) (bv-comp P1_P1_P3_HOLD  0b1)) (bv-and (bv-comp P1_P1_P3_READY_n  0b1) (bv-comp P1_P1_P3_NA_n  0b0)))   0b1)) ;1382
                                    P1_P1_P3_State <= #1 3'sb111; $display(";A 1384");		//(= P1_P1_P3_State    0b111)) ;1384
                                end
                                else begin
                                    $display(";A 1383");		//(= (bv-and (bv-or (bv-comp P1_P1_P3_RequestPending  0b1) (bv-comp P1_P1_P3_HOLD  0b1)) (bv-and (bv-comp P1_P1_P3_READY_n  0b1) (bv-comp P1_P1_P3_NA_n  0b0)))   0b0)) ;1383
                                    if (((((P1_P1_P3_RequestPending == 1'b1) & (P1_P1_P3_HOLD == 1'b0)) & (P1_P1_P3_READY_n == 1'b1)) & (P1_P1_P3_NA_n == 1'b0))) begin
                                        $display(";A 1385");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P1_P3_RequestPending  0b1) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_READY_n  0b1)) (bv-comp P1_P1_P3_NA_n  0b0))   0b1)) ;1385
                                        P1_P1_P3_State <= #1 3'sb110; $display(";A 1387");		//(= P1_P1_P3_State    0b110)) ;1387
                                    end
                                    else begin
                                        $display(";A 1386");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P1_P3_RequestPending  0b1) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_READY_n  0b1)) (bv-comp P1_P1_P3_NA_n  0b0))   0b0)) ;1386
                                        if ((((P1_P1_P3_RequestPending == 1'b0) & (P1_P1_P3_HOLD == 1'b0)) & (P1_P1_P3_READY_n == 1'b0))) begin
                                            $display(";A 1388");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_RequestPending  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_READY_n  0b0))   0b1)) ;1388
                                            P1_P1_P3_State <= #1 3'sb001; $display(";A 1390");		//(= P1_P1_P3_State    0b001)) ;1390
                                        end
                                        else begin
                                            $display(";A 1389");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_RequestPending  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_READY_n  0b0))   0b0)) ;1389
                                            if (((P1_P1_P3_HOLD == 1'b1) & (P1_P1_P3_READY_n == 1'b1))) begin
                                                $display(";A 1391");		//(= (bv-and (bv-comp P1_P1_P3_HOLD  0b1) (bv-comp P1_P1_P3_READY_n  0b1))   0b1)) ;1391
                                                P1_P1_P3_State <= #1 3'sb101; $display(";A 1393");		//(= P1_P1_P3_State    0b101)) ;1393
                                            end
                                            else begin
                                                $display(";A 1392");		//(= (bv-and (bv-comp P1_P1_P3_HOLD  0b1) (bv-comp P1_P1_P3_READY_n  0b1))   0b0)) ;1392
                                                P1_P1_P3_State <= #1 3'sb011; $display(";A 1394");		//(= P1_P1_P3_State    0b011)) ;1394
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P1_P1_P3_StateBS16 <= #1 P1_P1_P3_BS16_n; $display(";A 1395");		//(= P1_P1_P3_StateBS16    P1_P1_P3_BS16_n )) ;1395
                        if ((P1_P1_P3_BS16_n == 1'b0)) begin
                            $display(";A 1396");		//(= (bv-comp P1_P1_P3_BS16_n  0b0)   0b1)) ;1396
                            P1_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 1398");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000001)) ;1398
                        end
                        else begin
                            $display(";A 1397");		//(= (bv-comp P1_P1_P3_BS16_n  0b0)   0b0)) ;1397
                            P1_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 1399");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;1399
                        end
                        P1_P1_P3_StateNA <= #1 P1_P1_P3_NA_n; $display(";A 1400");		//(= P1_P1_P3_StateNA    P1_P1_P3_NA_n )) ;1400
                        P1_P1_P3_ADS_n <= #1 1'b1; $display(";A 1401");		//(= P1_P1_P3_ADS_n    0b1)) ;1401
                    end
                3'b100 :
                    begin
                        $display(";A 1402");		//(= P1_P1_P3_State    0b100)) ;1402
                        if ((((P1_P1_P3_NA_n == 1'b0) & (P1_P1_P3_HOLD == 1'b0)) & (P1_P1_P3_RequestPending == 1'b1))) begin
                            $display(";A 1403");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_NA_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b1))   0b1)) ;1403
                            P1_P1_P3_State <= #1 3'sb110; $display(";A 1405");		//(= P1_P1_P3_State    0b110)) ;1405
                        end
                        else begin
                            $display(";A 1404");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_NA_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b1))   0b0)) ;1404
                            if (((P1_P1_P3_NA_n == 1'b0) & ((P1_P1_P3_HOLD == 1'b1) | (P1_P1_P3_RequestPending == 1'b0)))) begin
                                $display(";A 1406");		//(= (bv-and (bv-comp P1_P1_P3_NA_n  0b0) (bv-or (bv-comp P1_P1_P3_HOLD  0b1) (bv-comp P1_P1_P3_RequestPending  0b0)))   0b1)) ;1406
                                P1_P1_P3_State <= #1 3'sb111; $display(";A 1408");		//(= P1_P1_P3_State    0b111)) ;1408
                            end
                            else begin
                                $display(";A 1407");		//(= (bv-and (bv-comp P1_P1_P3_NA_n  0b0) (bv-or (bv-comp P1_P1_P3_HOLD  0b1) (bv-comp P1_P1_P3_RequestPending  0b0)))   0b0)) ;1407
                                if ((P1_P1_P3_NA_n == 1'b1)) begin
                                    $display(";A 1409");		//(= (bv-comp P1_P1_P3_NA_n  0b1)   0b1)) ;1409
                                    P1_P1_P3_State <= #1 3'sb011; $display(";A 1411");		//(= P1_P1_P3_State    0b011)) ;1411
                                end
                                else begin
                                    $display(";A 1410");		//(= (bv-comp P1_P1_P3_NA_n  0b1)   0b0)) ;1410
                                    P1_P1_P3_State <= #1 3'sb100; $display(";A 1412");		//(= P1_P1_P3_State    0b100)) ;1412
                                end
                            end
                        end
                        P1_P1_P3_StateBS16 <= #1 P1_P1_P3_BS16_n; $display(";A 1413");		//(= P1_P1_P3_StateBS16    P1_P1_P3_BS16_n )) ;1413
                        if ((P1_P1_P3_BS16_n == 1'b0)) begin
                            $display(";A 1414");		//(= (bv-comp P1_P1_P3_BS16_n  0b0)   0b1)) ;1414
                            P1_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 1416");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000001)) ;1416
                        end
                        else begin
                            $display(";A 1415");		//(= (bv-comp P1_P1_P3_BS16_n  0b0)   0b0)) ;1415
                            P1_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 1417");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;1417
                        end
                        P1_P1_P3_StateNA <= #1 P1_P1_P3_NA_n; $display(";A 1418");		//(= P1_P1_P3_StateNA    P1_P1_P3_NA_n )) ;1418
                        P1_P1_P3_ADS_n <= #1 1'b1; $display(";A 1419");		//(= P1_P1_P3_ADS_n    0b1)) ;1419
                    end
                3'b101 :
                    begin
                        $display(";A 1420");		//(= P1_P1_P3_State    0b101)) ;1420
                        if (((P1_P1_P3_HOLD == 1'b0) & (P1_P1_P3_RequestPending == 1'b1))) begin
                            $display(";A 1421");		//(= (bv-and (bv-comp P1_P1_P3_HOLD  0b0) (bv-comp P1_P1_P3_RequestPending  0b1))   0b1)) ;1421
                            P1_P1_P3_State <= #1 3'sb010; $display(";A 1423");		//(= P1_P1_P3_State    0b010)) ;1423
                        end
                        else begin
                            $display(";A 1422");		//(= (bv-and (bv-comp P1_P1_P3_HOLD  0b0) (bv-comp P1_P1_P3_RequestPending  0b1))   0b0)) ;1422
                            if (((P1_P1_P3_HOLD == 1'b0) & (P1_P1_P3_RequestPending == 1'b0))) begin
                                $display(";A 1424");		//(= (bv-and (bv-comp P1_P1_P3_HOLD  0b0) (bv-comp P1_P1_P3_RequestPending  0b0))   0b1)) ;1424
                                P1_P1_P3_State <= #1 3'sb001; $display(";A 1426");		//(= P1_P1_P3_State    0b001)) ;1426
                            end
                            else begin
                                $display(";A 1425");		//(= (bv-and (bv-comp P1_P1_P3_HOLD  0b0) (bv-comp P1_P1_P3_RequestPending  0b0))   0b0)) ;1425
                                P1_P1_P3_State <= #1 3'sb101; $display(";A 1427");		//(= P1_P1_P3_State    0b101)) ;1427
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 1428");		//(= P1_P1_P3_State    0b110)) ;1428
                        P1_P1_P3_Address <= #1 ((P1_P1_P3_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 1429");		//(= P1_P1_P3_Address    (bv-smod (bv-sdiv P1_P1_P3_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;1429
                        P1_P1_P3_BE_n <= #1 P1_P1_P3_ByteEnable; $display(";A 1430");		//(= P1_P1_P3_BE_n    P1_P1_P3_ByteEnable )) ;1430
                        P1_P1_P3_M_IO_n <= #1 P1_P1_P3_MemoryFetch; $display(";A 1431");		//(= P1_P1_P3_M_IO_n    P1_P1_P3_MemoryFetch )) ;1431
                        if ((P1_P1_P3_ReadRequest == 1'b1)) begin
                            $display(";A 1432");		//(= (bv-comp P1_P1_P3_ReadRequest  0b1)   0b1)) ;1432
                            P1_P1_P3_W_R_n <= #1 1'b0; $display(";A 1434");		//(= P1_P1_P3_W_R_n    0b0)) ;1434
                        end
                        else begin
                            $display(";A 1433");		//(= (bv-comp P1_P1_P3_ReadRequest  0b1)   0b0)) ;1433
                            P1_P1_P3_W_R_n <= #1 1'b1; $display(";A 1435");		//(= P1_P1_P3_W_R_n    0b1)) ;1435
                        end
                        if ((P1_P1_P3_CodeFetch == 1'b1)) begin
                            $display(";A 1436");		//(= (bv-comp P1_P1_P3_CodeFetch  0b1)   0b1)) ;1436
                            P1_P1_P3_D_C_n <= #1 1'b0; $display(";A 1438");		//(= P1_P1_P3_D_C_n    0b0)) ;1438
                        end
                        else begin
                            $display(";A 1437");		//(= (bv-comp P1_P1_P3_CodeFetch  0b1)   0b0)) ;1437
                            P1_P1_P3_D_C_n <= #1 1'b1; $display(";A 1439");		//(= P1_P1_P3_D_C_n    0b1)) ;1439
                        end
                        P1_P1_P3_ADS_n <= #1 1'b0; $display(";A 1440");		//(= P1_P1_P3_ADS_n    0b0)) ;1440
                        if ((P1_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 1441");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1441
                            P1_P1_P3_State <= #1 3'sb100; $display(";A 1443");		//(= P1_P1_P3_State    0b100)) ;1443
                        end
                        else begin
                            $display(";A 1442");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1442
                            P1_P1_P3_State <= #1 3'sb110; $display(";A 1444");		//(= P1_P1_P3_State    0b110)) ;1444
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 1445");		//(= P1_P1_P3_State    0b111)) ;1445
                        if ((((P1_P1_P3_READY_n == 1'b1) & (P1_P1_P3_RequestPending == 1'b1)) & (P1_P1_P3_HOLD == 1'b0))) begin
                            $display(";A 1446");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b1) (bv-comp P1_P1_P3_RequestPending  0b1)) (bv-comp P1_P1_P3_HOLD  0b0))   0b1)) ;1446
                            P1_P1_P3_State <= #1 3'sb110; $display(";A 1448");		//(= P1_P1_P3_State    0b110)) ;1448
                        end
                        else begin
                            $display(";A 1447");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b1) (bv-comp P1_P1_P3_RequestPending  0b1)) (bv-comp P1_P1_P3_HOLD  0b0))   0b0)) ;1447
                            if (((P1_P1_P3_READY_n == 1'b0) & (P1_P1_P3_HOLD == 1'b1))) begin
                                $display(";A 1449");		//(= (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b1))   0b1)) ;1449
                                P1_P1_P3_State <= #1 3'sb101; $display(";A 1451");		//(= P1_P1_P3_State    0b101)) ;1451
                            end
                            else begin
                                $display(";A 1450");		//(= (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b1))   0b0)) ;1450
                                if ((((P1_P1_P3_READY_n == 1'b0) & (P1_P1_P3_HOLD == 1'b0)) & (P1_P1_P3_RequestPending == 1'b1))) begin
                                    $display(";A 1452");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b1))   0b1)) ;1452
                                    P1_P1_P3_State <= #1 3'sb010; $display(";A 1454");		//(= P1_P1_P3_State    0b010)) ;1454
                                end
                                else begin
                                    $display(";A 1453");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b1))   0b0)) ;1453
                                    if ((((P1_P1_P3_READY_n == 1'b0) & (P1_P1_P3_HOLD == 1'b0)) & (P1_P1_P3_RequestPending == 1'b0))) begin
                                        $display(";A 1455");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b0))   0b1)) ;1455
                                        P1_P1_P3_State <= #1 3'sb001; $display(";A 1457");		//(= P1_P1_P3_State    0b001)) ;1457
                                    end
                                    else begin
                                        $display(";A 1456");		//(= (bv-and (bv-and (bv-comp P1_P1_P3_READY_n  0b0) (bv-comp P1_P1_P3_HOLD  0b0)) (bv-comp P1_P1_P3_RequestPending  0b0))   0b0)) ;1456
                                        P1_P1_P3_State <= #1 3'sb111; $display(";A 1458");		//(= P1_P1_P3_State    0b111)) ;1458
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2030
    always @(posedge P1_P1_P3_RESET or posedge P1_P1_P3_CLOCK) begin
        if ((P1_P1_P3_RESET == 1'b1)) begin
            $display(";A 1459");		//(= (bv-comp P1_P1_P3_RESET  0b1)   0b1)) ;1459
            P1_P1_P3_State2 = 4'sb0000; $display(";A 1461");		//(= P1_P1_P3_State2    0b0000)) ;1461
            P1_P1_P3_InstQueue[0] = 8'b00000000; $display(";A 1462");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1462
            P1_P1_P3_InstQueue[1] = 8'b00000000; $display(";A 1463");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1463
            P1_P1_P3_InstQueue[2] = 8'b00000000; $display(";A 1464");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1464
            P1_P1_P3_InstQueue[3] = 8'b00000000; $display(";A 1465");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1465
            P1_P1_P3_InstQueue[4] = 8'b00000000; $display(";A 1466");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1466
            P1_P1_P3_InstQueue[5] = 8'b00000000; $display(";A 1467");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1467
            P1_P1_P3_InstQueue[6] = 8'b00000000; $display(";A 1468");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1468
            P1_P1_P3_InstQueue[7] = 8'b00000000; $display(";A 1469");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1469
            P1_P1_P3_InstQueue[8] = 8'b00000000; $display(";A 1470");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1470
            P1_P1_P3_InstQueue[9] = 8'b00000000; $display(";A 1471");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1471
            P1_P1_P3_InstQueue[10] = 8'b00000000; $display(";A 1472");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1472
            P1_P1_P3_InstQueue[11] = 8'b00000000; $display(";A 1473");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1473
            P1_P1_P3_InstQueue[12] = 8'b00000000; $display(";A 1474");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1474
            P1_P1_P3_InstQueue[13] = 8'b00000000; $display(";A 1475");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1475
            P1_P1_P3_InstQueue[14] = 8'b00000000; $display(";A 1476");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1476
            P1_P1_P3_InstQueue[15] = 8'b00000000; $display(";A 1477");		//(= P1_P1_P3_InstQueue    0b00000000)) ;1477
            P1_P1_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 1478");		//(= P1_P1_P3_InstQueueRd_Addr    0b00000)) ;1478
            P1_P1_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 1479");		//(= P1_P1_P3_InstQueueWr_Addr    0b00000)) ;1479
            P1_P1_P3_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 1480");		//(= P1_P1_P3_InstAddrPointer    0b00000000000000000000000000000000)) ;1480
            P1_P1_P3_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 1481");		//(= P1_P1_P3_PhyAddrPointer    0b00000000000000000000000000000000)) ;1481
            P1_P1_P3_Extended = 1'b0; $display(";A 1482");		//(= P1_P1_P3_Extended    0b0)) ;1482
            P1_P1_P3_More = 1'b0; $display(";A 1483");		//(= P1_P1_P3_More    0b0)) ;1483
            P1_P1_P3_Flush = 1'b0; $display(";A 1484");		//(= P1_P1_P3_Flush    0b0)) ;1484
            P1_P1_P3_lWord = 16'sb0000000000000000; $display(";A 1485");		//(= P1_P1_P3_lWord    0b0000000000000000)) ;1485
            P1_P1_P3_uWord = 15'sb000000000000000; $display(";A 1486");		//(= P1_P1_P3_uWord    0b000000000000000)) ;1486
            P1_P1_P3_fWord = 32'sb00000000000000000000000000000000; $display(";A 1487");		//(= P1_P1_P3_fWord    0b00000000000000000000000000000000)) ;1487
            P1_P1_P3_CodeFetch <= #1 1'b0; $display(";A 1488");		//(= P1_P1_P3_CodeFetch    0b0)) ;1488
            P1_P1_P3_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 1489");		//(= P1_P1_P3_Datao    0b00000000000000000000000000000000)) ;1489
            P1_P1_P3_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 1490");		//(= P1_P1_P3_EAX    0b00000000000000000000000000000000)) ;1490
            P1_P1_P3_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 1491");		//(= P1_P1_P3_EBX    0b00000000000000000000000000000000)) ;1491
            P1_P1_P3_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 1492");		//(= P1_P1_P3_rEIP    0b00000000000000000000000000000000)) ;1492
            P1_P1_P3_ReadRequest <= #1 1'b0; $display(";A 1493");		//(= P1_P1_P3_ReadRequest    0b0)) ;1493
            P1_P1_P3_MemoryFetch <= #1 1'b0; $display(";A 1494");		//(= P1_P1_P3_MemoryFetch    0b0)) ;1494
            P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1495");		//(= P1_P1_P3_RequestPending    0b0)) ;1495
        end
        else begin
            $display(";A 1460");		//(= (bv-comp P1_P1_P3_RESET  0b1)   0b0)) ;1460
            case (P1_P1_P3_State2)
                4'b0000 :
                    begin
                        $display(";A 1496");		//(= P1_P1_P3_State2    0b0000)) ;1496
                        P1_P1_P3_PhyAddrPointer = P1_P1_P3_rEIP; $display(";A 1497");		//(= P1_P1_P3_PhyAddrPointer    P1_P1_P3_rEIP )) ;1497
                        P1_P1_P3_InstAddrPointer = P1_P1_P3_PhyAddrPointer; $display(";A 1498");		//(= P1_P1_P3_InstAddrPointer    P1_P1_P3_PhyAddrPointer )) ;1498
                        P1_P1_P3_State2 = 4'sb0001; $display(";A 1499");		//(= P1_P1_P3_State2    0b0001)) ;1499
                        P1_P1_P3_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 1500");		//(= P1_P1_P3_rEIP    0b00000000000011111111111111110000)) ;1500
                        P1_P1_P3_ReadRequest <= #1 1'b1; $display(";A 1501");		//(= P1_P1_P3_ReadRequest    0b1)) ;1501
                        P1_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 1502");		//(= P1_P1_P3_MemoryFetch    0b1)) ;1502
                        P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1503");		//(= P1_P1_P3_RequestPending    0b1)) ;1503
                    end
                4'b0001 :
                    begin
                        $display(";A 1504");		//(= P1_P1_P3_State2    0b0001)) ;1504
                        P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1505");		//(= P1_P1_P3_RequestPending    0b1)) ;1505
                        P1_P1_P3_ReadRequest <= #1 1'b1; $display(";A 1506");		//(= P1_P1_P3_ReadRequest    0b1)) ;1506
                        P1_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 1507");		//(= P1_P1_P3_MemoryFetch    0b1)) ;1507
                        P1_P1_P3_CodeFetch <= #1 1'b1; $display(";A 1508");		//(= P1_P1_P3_CodeFetch    0b1)) ;1508
                        if ((P1_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 1509");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1509
                            P1_P1_P3_State2 = 4'sb0010; $display(";A 1511");		//(= P1_P1_P3_State2    0b0010)) ;1511
                        end
                        else begin
                            $display(";A 1510");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1510
                            P1_P1_P3_State2 = 4'sb0001; $display(";A 1512");		//(= P1_P1_P3_State2    0b0001)) ;1512
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 1513");		//(= P1_P1_P3_State2    0b0010)) ;1513
                        P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1514");		//(= P1_P1_P3_RequestPending    0b0)) ;1514
                        P1_P1_P3_InstQueue[P1_P1_P3_InstQueueWr_Addr] = (P1_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 1515");		//(= P1_P1_P3_InstQueue    (bv-smod P1_P1_P3_Datai  0b00000000000000000000000100000000))) ;1515
                        P1_P1_P3_InstQueueWr_Addr = ((P1_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1516");		//(= P1_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1516
                        P1_P1_P3_InstQueue[P1_P1_P3_InstQueueWr_Addr] = (P1_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 1517");		//(= P1_P1_P3_InstQueue    (bv-smod P1_P1_P3_Datai  0b00000000000000000000000100000000))) ;1517
                        P1_P1_P3_InstQueueWr_Addr = ((P1_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1518");		//(= P1_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1518
                        if ((P1_P1_P3_StateBS16 == 1'b1)) begin
                            $display(";A 1519");		//(= (bv-comp P1_P1_P3_StateBS16  0b1)   0b1)) ;1519
                            P1_P1_P3_InstQueue[P1_P1_P3_InstQueueWr_Addr] = ((P1_P1_P3_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 1521");		//(= P1_P1_P3_InstQueue    (bv-smod (bv-sdiv P1_P1_P3_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;1521
                            P1_P1_P3_InstQueueWr_Addr = ((P1_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1522");		//(= P1_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1522
                            P1_P1_P3_InstQueue[P1_P1_P3_InstQueueWr_Addr] = ((P1_P1_P3_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 1523");		//(= P1_P1_P3_InstQueue    (bv-smod (bv-sdiv P1_P1_P3_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;1523
                            P1_P1_P3_InstQueueWr_Addr = ((P1_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1524");		//(= P1_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1524
                            P1_P1_P3_PhyAddrPointer = (P1_P1_P3_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 1525");		//(= P1_P1_P3_PhyAddrPointer    (bv-add P1_P1_P3_PhyAddrPointer  0b00000000000000000000000000000100))) ;1525
                            P1_P1_P3_State2 = 4'sb0101; $display(";A 1526");		//(= P1_P1_P3_State2    0b0101)) ;1526
                        end
                        else begin
                            $display(";A 1520");		//(= (bv-comp P1_P1_P3_StateBS16  0b1)   0b0)) ;1520
                            P1_P1_P3_PhyAddrPointer = (P1_P1_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1527");		//(= P1_P1_P3_PhyAddrPointer    (bv-add P1_P1_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;1527
                            if ((P1_P1_P3_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 1528");		//(= (bool-to-bv (bv-slt P1_P1_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;1528
                                P1_P1_P3_rEIP <= #1 (-P1_P1_P3_PhyAddrPointer); $display(";A 1530");		//(= P1_P1_P3_rEIP    (bv-neg P1_P1_P3_PhyAddrPointer ))) ;1530
                            end
                            else begin
                                $display(";A 1529");		//(= (bool-to-bv (bv-slt P1_P1_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;1529
                                P1_P1_P3_rEIP <= #1 P1_P1_P3_PhyAddrPointer; $display(";A 1531");		//(= P1_P1_P3_rEIP    P1_P1_P3_PhyAddrPointer )) ;1531
                            end
                            P1_P1_P3_State2 = 4'sb0011; $display(";A 1532");		//(= P1_P1_P3_State2    0b0011)) ;1532
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 1533");		//(= P1_P1_P3_State2    0b0011)) ;1533
                        P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1534");		//(= P1_P1_P3_RequestPending    0b1)) ;1534
                        if ((P1_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 1535");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1535
                            P1_P1_P3_State2 = 4'sb0100; $display(";A 1537");		//(= P1_P1_P3_State2    0b0100)) ;1537
                        end
                        else begin
                            $display(";A 1536");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1536
                            P1_P1_P3_State2 = 4'sb0011; $display(";A 1538");		//(= P1_P1_P3_State2    0b0011)) ;1538
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 1539");		//(= P1_P1_P3_State2    0b0100)) ;1539
                        P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1540");		//(= P1_P1_P3_RequestPending    0b0)) ;1540
                        P1_P1_P3_InstQueue[P1_P1_P3_InstQueueWr_Addr] = (P1_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 1541");		//(= P1_P1_P3_InstQueue    (bv-smod P1_P1_P3_Datai  0b00000000000000000000000100000000))) ;1541
                        P1_P1_P3_InstQueueWr_Addr = ((P1_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1542");		//(= P1_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1542
                        P1_P1_P3_InstQueue[P1_P1_P3_InstQueueWr_Addr] = (P1_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 1543");		//(= P1_P1_P3_InstQueue    (bv-smod P1_P1_P3_Datai  0b00000000000000000000000100000000))) ;1543
                        P1_P1_P3_InstQueueWr_Addr = ((P1_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1544");		//(= P1_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1544
                        P1_P1_P3_PhyAddrPointer = (P1_P1_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1545");		//(= P1_P1_P3_PhyAddrPointer    (bv-add P1_P1_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;1545
                        P1_P1_P3_State2 = 4'sb0101; $display(";A 1546");		//(= P1_P1_P3_State2    0b0101)) ;1546
                    end
                4'b0101 :
                    begin
                        $display(";A 1547");		//(= P1_P1_P3_State2    0b0101)) ;1547
                        case (P1_P1_P3_InstQueue[P1_P1_P3_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 1548");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b10010000)) ;1548
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1549");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1549
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1550");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1550
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1551");		//(= P1_P1_P3_Flush    0b0)) ;1551
                                    P1_P1_P3_More = 1'b0; $display(";A 1552");		//(= P1_P1_P3_More    0b0)) ;1552
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 1553");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b01100110)) ;1553
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1554");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1554
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1555");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1555
                                    P1_P1_P3_Extended = 1'b1; $display(";A 1556");		//(= P1_P1_P3_Extended    0b1)) ;1556
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1557");		//(= P1_P1_P3_Flush    0b0)) ;1557
                                    P1_P1_P3_More = 1'b0; $display(";A 1558");		//(= P1_P1_P3_More    0b0)) ;1558
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 1559");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b11101011)) ;1559
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 1560");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;1560
                                        if ((P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 1562");		//(= (bool-to-bv (bv-gt P1_P1_P3_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;1562
                                            P1_P1_P3_PhyAddrPointer = ((P1_P1_P3_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 1564");		//(= P1_P1_P3_PhyAddrPointer    (bv-sub (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P1_P1_P3_InstQueue 0 )))) ;1564
                                            P1_P1_P3_InstAddrPointer = P1_P1_P3_PhyAddrPointer; $display(";A 1565");		//(= P1_P1_P3_InstAddrPointer    P1_P1_P3_PhyAddrPointer )) ;1565
                                        end
                                        else begin
                                            $display(";A 1563");		//(= (bool-to-bv (bv-gt P1_P1_P3_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;1563
                                            P1_P1_P3_PhyAddrPointer = ((P1_P1_P3_InstAddrPointer + 32'b00000000000000000000000000000010) + P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 1566");		//(= P1_P1_P3_PhyAddrPointer    (bv-add (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000010) P1_P1_P3_InstQueue 0 ))) ;1566
                                            P1_P1_P3_InstAddrPointer = P1_P1_P3_PhyAddrPointer; $display(";A 1567");		//(= P1_P1_P3_InstAddrPointer    P1_P1_P3_PhyAddrPointer )) ;1567
                                        end
                                        P1_P1_P3_Flush = 1'b1; $display(";A 1568");		//(= P1_P1_P3_Flush    0b1)) ;1568
                                        P1_P1_P3_More = 1'b0; $display(";A 1569");		//(= P1_P1_P3_More    0b0)) ;1569
                                    end
                                    else begin
                                        $display(";A 1561");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;1561
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1570");		//(= P1_P1_P3_Flush    0b0)) ;1570
                                        P1_P1_P3_More = 1'b1; $display(";A 1571");		//(= P1_P1_P3_More    0b1)) ;1571
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 1572");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b11101001)) ;1572
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 1573");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;1573
                                        P1_P1_P3_PhyAddrPointer = ((P1_P1_P3_InstAddrPointer + 32'b00000000000000000000000000000101) + P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 1575");		//(= P1_P1_P3_PhyAddrPointer    (bv-add (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000101) P1_P1_P3_InstQueue 0 ))) ;1575
                                        P1_P1_P3_InstAddrPointer = P1_P1_P3_PhyAddrPointer; $display(";A 1576");		//(= P1_P1_P3_InstAddrPointer    P1_P1_P3_PhyAddrPointer )) ;1576
                                        P1_P1_P3_Flush = 1'b1; $display(";A 1577");		//(= P1_P1_P3_Flush    0b1)) ;1577
                                        P1_P1_P3_More = 1'b0; $display(";A 1578");		//(= P1_P1_P3_More    0b0)) ;1578
                                    end
                                    else begin
                                        $display(";A 1574");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;1574
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1579");		//(= P1_P1_P3_Flush    0b0)) ;1579
                                        P1_P1_P3_More = 1'b1; $display(";A 1580");		//(= P1_P1_P3_More    0b1)) ;1580
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 1581");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b11101010)) ;1581
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1582");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1582
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1583");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1583
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1584");		//(= P1_P1_P3_Flush    0b0)) ;1584
                                    P1_P1_P3_More = 1'b0; $display(";A 1585");		//(= P1_P1_P3_More    0b0)) ;1585
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 1586");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b10110000)) ;1586
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1587");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1587
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1588");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1588
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1589");		//(= P1_P1_P3_Flush    0b0)) ;1589
                                    P1_P1_P3_More = 1'b0; $display(";A 1590");		//(= P1_P1_P3_More    0b0)) ;1590
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 1591");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b10111000)) ;1591
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 1592");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;1592
                                        P1_P1_P3_EAX <= #1 ((((P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 1594");		//(= P1_P1_P3_EAX    (bv-add (bv-add (bv-add (bv-mul P1_P1_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P1_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P1_P3_InstQueue 0  0b00000000000000000000000100000000)) P1_P1_P3_InstQueue 0 ))) ;1594
                                        P1_P1_P3_More = 1'b0; $display(";A 1595");		//(= P1_P1_P3_More    0b0)) ;1595
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1596");		//(= P1_P1_P3_Flush    0b0)) ;1596
                                        P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 1597");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;1597
                                        P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 1598");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;1598
                                    end
                                    else begin
                                        $display(";A 1593");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;1593
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1599");		//(= P1_P1_P3_Flush    0b0)) ;1599
                                        P1_P1_P3_More = 1'b1; $display(";A 1600");		//(= P1_P1_P3_More    0b1)) ;1600
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 1601");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b10111011)) ;1601
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 1602");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;1602
                                        P1_P1_P3_EBX <= #1 ((((P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P1_P3_InstQueue[((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 1604");		//(= P1_P1_P3_EBX    (bv-add (bv-add (bv-add (bv-mul P1_P1_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P1_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P1_P3_InstQueue 0  0b00000000000000000000000100000000)) P1_P1_P3_InstQueue 0 ))) ;1604
                                        P1_P1_P3_More = 1'b0; $display(";A 1605");		//(= P1_P1_P3_More    0b0)) ;1605
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1606");		//(= P1_P1_P3_Flush    0b0)) ;1606
                                        P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 1607");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;1607
                                        P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 1608");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;1608
                                    end
                                    else begin
                                        $display(";A 1603");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;1603
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1609");		//(= P1_P1_P3_Flush    0b0)) ;1609
                                        P1_P1_P3_More = 1'b1; $display(";A 1610");		//(= P1_P1_P3_More    0b1)) ;1610
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 1611");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b10001011)) ;1611
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1612");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1612
                                        if ((P1_P1_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 1614");		//(= (bool-to-bv (bv-slt P1_P1_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;1614
                                            P1_P1_P3_rEIP <= #1 (-P1_P1_P3_EBX); $display(";A 1616");		//(= P1_P1_P3_rEIP    (bv-neg P1_P1_P3_EBX ))) ;1616
                                        end
                                        else begin
                                            $display(";A 1615");		//(= (bool-to-bv (bv-slt P1_P1_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;1615
                                            P1_P1_P3_rEIP <= #1 P1_P1_P3_EBX; $display(";A 1617");		//(= P1_P1_P3_rEIP    P1_P1_P3_EBX )) ;1617
                                        end
                                        P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1618");		//(= P1_P1_P3_RequestPending    0b1)) ;1618
                                        P1_P1_P3_ReadRequest <= #1 1'b1; $display(";A 1619");		//(= P1_P1_P3_ReadRequest    0b1)) ;1619
                                        P1_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 1620");		//(= P1_P1_P3_MemoryFetch    0b1)) ;1620
                                        P1_P1_P3_CodeFetch <= #1 1'b0; $display(";A 1621");		//(= P1_P1_P3_CodeFetch    0b0)) ;1621
                                        if ((P1_P1_P3_READY_n == 1'b0)) begin
                                            $display(";A 1622");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1622
                                            P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1624");		//(= P1_P1_P3_RequestPending    0b0)) ;1624
                                            P1_P1_P3_uWord = (P1_P1_P3_Datai % 32'b00000000000000001000000000000000); $display(";A 1625");		//(= P1_P1_P3_uWord    (bv-smod P1_P1_P3_Datai  0b00000000000000001000000000000000))) ;1625
                                            if ((P1_P1_P3_StateBS16 == 1'b1)) begin
                                                $display(";A 1626");		//(= (bv-comp P1_P1_P3_StateBS16  0b1)   0b1)) ;1626
                                                P1_P1_P3_lWord = (P1_P1_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 1628");		//(= P1_P1_P3_lWord    (bv-smod P1_P1_P3_Datai  0b00000000000000010000000000000000))) ;1628
                                            end
                                            else begin
                                                $display(";A 1627");		//(= (bv-comp P1_P1_P3_StateBS16  0b1)   0b0)) ;1627
                                                P1_P1_P3_rEIP <= #1 (P1_P1_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 1629");		//(= P1_P1_P3_rEIP    (bv-add P1_P1_P3_rEIP  0b00000000000000000000000000000010))) ;1629
                                                P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1630");		//(= P1_P1_P3_RequestPending    0b1)) ;1630
                                                if ((P1_P1_P3_READY_n == 1'b0)) begin
                                                    $display(";A 1631");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1631
                                                    P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1633");		//(= P1_P1_P3_RequestPending    0b0)) ;1633
                                                    P1_P1_P3_lWord = (P1_P1_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 1634");		//(= P1_P1_P3_lWord    (bv-smod P1_P1_P3_Datai  0b00000000000000010000000000000000))) ;1634
                                                end
                                                else begin
                                                    $display(";A 1632");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1632
                                                end
                                            end
                                            if ((P1_P1_P3_READY_n == 1'b0)) begin
                                                $display(";A 1635");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1635
                                                P1_P1_P3_EAX <= #1 ((P1_P1_P3_uWord * 32'b00000000000000010000000000000000) + P1_P1_P3_lWord); $display(";A 1637");		//(= P1_P1_P3_EAX    (bv-add (bv-mul P1_P1_P3_uWord  0b00000000000000010000000000000000) P1_P1_P3_lWord ))) ;1637
                                                P1_P1_P3_More = 1'b0; $display(";A 1638");		//(= P1_P1_P3_More    0b0)) ;1638
                                                P1_P1_P3_Flush = 1'b0; $display(";A 1639");		//(= P1_P1_P3_Flush    0b0)) ;1639
                                                P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1640");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;1640
                                                P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1641");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1641
                                            end
                                            else begin
                                                $display(";A 1636");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1636
                                            end
                                        end
                                        else begin
                                            $display(";A 1623");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1623
                                        end
                                    end
                                    else begin
                                        $display(";A 1613");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1613
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1642");		//(= P1_P1_P3_Flush    0b0)) ;1642
                                        P1_P1_P3_More = 1'b1; $display(";A 1643");		//(= P1_P1_P3_More    0b1)) ;1643
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 1644");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b10001001)) ;1644
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1645");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1645
                                        if ((P1_P1_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 1647");		//(= (bool-to-bv (bv-slt P1_P1_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;1647
                                            P1_P1_P3_rEIP <= #1 P1_P1_P3_EBX; $display(";A 1649");		//(= P1_P1_P3_rEIP    P1_P1_P3_EBX )) ;1649
                                        end
                                        else begin
                                            $display(";A 1648");		//(= (bool-to-bv (bv-slt P1_P1_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;1648
                                            P1_P1_P3_rEIP <= #1 P1_P1_P3_EBX; $display(";A 1650");		//(= P1_P1_P3_rEIP    P1_P1_P3_EBX )) ;1650
                                        end
                                        P1_P1_P3_lWord = (P1_P1_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 1651");		//(= P1_P1_P3_lWord    (bv-smod P1_P1_P3_EAX  0b00000000000000010000000000000000))) ;1651
                                        P1_P1_P3_uWord = ((P1_P1_P3_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 1652");		//(= P1_P1_P3_uWord    (bv-smod (bv-sdiv P1_P1_P3_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;1652
                                        P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1653");		//(= P1_P1_P3_RequestPending    0b1)) ;1653
                                        P1_P1_P3_ReadRequest <= #1 1'b0; $display(";A 1654");		//(= P1_P1_P3_ReadRequest    0b0)) ;1654
                                        P1_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 1655");		//(= P1_P1_P3_MemoryFetch    0b1)) ;1655
                                        P1_P1_P3_CodeFetch <= #1 1'b0; $display(";A 1656");		//(= P1_P1_P3_CodeFetch    0b0)) ;1656
                                        if (((P1_P1_P3_State == 32'b00000000000000000000000000000010) | (P1_P1_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 1657");		//(= (bv-or (bv-comp P1_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P3_State  0b00000000000000000000000000000100))   0b1)) ;1657
                                            P1_P1_P3_Datao <= #1 ((P1_P1_P3_uWord * 32'b00000000000000010000000000000000) + P1_P1_P3_lWord); $display(";A 1659");		//(= P1_P1_P3_Datao    (bv-add (bv-mul P1_P1_P3_uWord  0b00000000000000010000000000000000) P1_P1_P3_lWord ))) ;1659
                                            if ((P1_P1_P3_READY_n == 1'b0)) begin
                                                $display(";A 1660");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1660
                                                P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1662");		//(= P1_P1_P3_RequestPending    0b0)) ;1662
                                                if ((P1_P1_P3_StateBS16 == 1'b0)) begin
                                                    $display(";A 1663");		//(= (bv-comp P1_P1_P3_StateBS16  0b0)   0b1)) ;1663
                                                    P1_P1_P3_rEIP <= #1 (P1_P1_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 1665");		//(= P1_P1_P3_rEIP    (bv-add P1_P1_P3_rEIP  0b00000000000000000000000000000010))) ;1665
                                                    P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1666");		//(= P1_P1_P3_RequestPending    0b1)) ;1666
                                                    P1_P1_P3_ReadRequest <= #1 1'b0; $display(";A 1667");		//(= P1_P1_P3_ReadRequest    0b0)) ;1667
                                                    P1_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 1668");		//(= P1_P1_P3_MemoryFetch    0b1)) ;1668
                                                    P1_P1_P3_CodeFetch <= #1 1'b0; $display(";A 1669");		//(= P1_P1_P3_CodeFetch    0b0)) ;1669
                                                    P1_P1_P3_State2 = 4'sb0110; $display(";A 1670");		//(= P1_P1_P3_State2    0b0110)) ;1670
                                                end
                                                else begin
                                                    $display(";A 1664");		//(= (bv-comp P1_P1_P3_StateBS16  0b0)   0b0)) ;1664
                                                end
                                                P1_P1_P3_More = 1'b0; $display(";A 1671");		//(= P1_P1_P3_More    0b0)) ;1671
                                                P1_P1_P3_Flush = 1'b0; $display(";A 1672");		//(= P1_P1_P3_Flush    0b0)) ;1672
                                                P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1673");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;1673
                                                P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1674");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1674
                                            end
                                            else begin
                                                $display(";A 1661");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1661
                                            end
                                        end
                                        else begin
                                            $display(";A 1658");		//(= (bv-or (bv-comp P1_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P3_State  0b00000000000000000000000000000100))   0b0)) ;1658
                                        end
                                    end
                                    else begin
                                        $display(";A 1646");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1646
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1675");		//(= P1_P1_P3_Flush    0b0)) ;1675
                                        P1_P1_P3_More = 1'b1; $display(";A 1676");		//(= P1_P1_P3_More    0b1)) ;1676
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 1677");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b11100100)) ;1677
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1678");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1678
                                        P1_P1_P3_rEIP <= #1 (P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 1680");		//(= P1_P1_P3_rEIP    (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;1680
                                        P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1681");		//(= P1_P1_P3_RequestPending    0b1)) ;1681
                                        P1_P1_P3_ReadRequest <= #1 1'b1; $display(";A 1682");		//(= P1_P1_P3_ReadRequest    0b1)) ;1682
                                        P1_P1_P3_MemoryFetch <= #1 1'b0; $display(";A 1683");		//(= P1_P1_P3_MemoryFetch    0b0)) ;1683
                                        P1_P1_P3_CodeFetch <= #1 1'b0; $display(";A 1684");		//(= P1_P1_P3_CodeFetch    0b0)) ;1684
                                        if ((P1_P1_P3_READY_n == 1'b0)) begin
                                            $display(";A 1685");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1685
                                            P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1687");		//(= P1_P1_P3_RequestPending    0b0)) ;1687
                                            P1_P1_P3_EAX <= #1 P1_P1_P3_Datai; $display(";A 1688");		//(= P1_P1_P3_EAX    P1_P1_P3_Datai )) ;1688
                                            P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1689");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;1689
                                            P1_P1_P3_InstQueueRd_Addr = (P1_P1_P3_InstQueueRd_Addr + 5'b00010); $display(";A 1690");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-add P1_P1_P3_InstQueueRd_Addr  0b00010))) ;1690
                                            P1_P1_P3_Flush = 1'b0; $display(";A 1691");		//(= P1_P1_P3_Flush    0b0)) ;1691
                                            P1_P1_P3_More = 1'b0; $display(";A 1692");		//(= P1_P1_P3_More    0b0)) ;1692
                                        end
                                        else begin
                                            $display(";A 1686");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1686
                                        end
                                    end
                                    else begin
                                        $display(";A 1679");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1679
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1693");		//(= P1_P1_P3_Flush    0b0)) ;1693
                                        P1_P1_P3_More = 1'b1; $display(";A 1694");		//(= P1_P1_P3_More    0b1)) ;1694
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 1695");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b11100110)) ;1695
                                    if (((P1_P1_P3_InstQueueWr_Addr - P1_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 1696");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;1696
                                        P1_P1_P3_rEIP <= #1 (P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 1698");		//(= P1_P1_P3_rEIP    (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;1698
                                        P1_P1_P3_RequestPending <= #1 1'b1; $display(";A 1699");		//(= P1_P1_P3_RequestPending    0b1)) ;1699
                                        P1_P1_P3_ReadRequest <= #1 1'b0; $display(";A 1700");		//(= P1_P1_P3_ReadRequest    0b0)) ;1700
                                        P1_P1_P3_MemoryFetch <= #1 1'b0; $display(";A 1701");		//(= P1_P1_P3_MemoryFetch    0b0)) ;1701
                                        P1_P1_P3_CodeFetch <= #1 1'b0; $display(";A 1702");		//(= P1_P1_P3_CodeFetch    0b0)) ;1702
                                        if (((P1_P1_P3_State == 32'b00000000000000000000000000000010) | (P1_P1_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 1703");		//(= (bv-or (bv-comp P1_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P3_State  0b00000000000000000000000000000100))   0b1)) ;1703
                                            P1_P1_P3_fWord = (P1_P1_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 1705");		//(= P1_P1_P3_fWord    (bv-smod P1_P1_P3_EAX  0b00000000000000010000000000000000))) ;1705
                                            P1_P1_P3_Datao <= #1 P1_P1_P3_fWord; $display(";A 1706");		//(= P1_P1_P3_Datao    P1_P1_P3_fWord )) ;1706
                                            if ((P1_P1_P3_READY_n == 1'b0)) begin
                                                $display(";A 1707");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1707
                                                P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1709");		//(= P1_P1_P3_RequestPending    0b0)) ;1709
                                                P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1710");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;1710
                                                P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1711");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1711
                                                P1_P1_P3_Flush = 1'b0; $display(";A 1712");		//(= P1_P1_P3_Flush    0b0)) ;1712
                                                P1_P1_P3_More = 1'b0; $display(";A 1713");		//(= P1_P1_P3_More    0b0)) ;1713
                                            end
                                            else begin
                                                $display(";A 1708");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1708
                                            end
                                        end
                                        else begin
                                            $display(";A 1704");		//(= (bv-or (bv-comp P1_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P1_P3_State  0b00000000000000000000000000000100))   0b0)) ;1704
                                        end
                                    end
                                    else begin
                                        $display(";A 1697");		//(= (bool-to-bv (bv-ge (bv-sub P1_P1_P3_InstQueueWr_Addr  P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;1697
                                        P1_P1_P3_Flush = 1'b0; $display(";A 1714");		//(= P1_P1_P3_Flush    0b0)) ;1714
                                        P1_P1_P3_More = 1'b1; $display(";A 1715");		//(= P1_P1_P3_More    0b1)) ;1715
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 1716");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b00000100)) ;1716
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1717");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1717
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1718");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1718
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1719");		//(= P1_P1_P3_Flush    0b0)) ;1719
                                    P1_P1_P3_More = 1'b0; $display(";A 1720");		//(= P1_P1_P3_More    0b0)) ;1720
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 1721");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b00000101)) ;1721
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1722");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1722
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1723");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1723
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1724");		//(= P1_P1_P3_Flush    0b0)) ;1724
                                    P1_P1_P3_More = 1'b0; $display(";A 1725");		//(= P1_P1_P3_More    0b0)) ;1725
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 1726");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b11010000)) ;1726
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1727");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;1727
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1728");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1728
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1729");		//(= P1_P1_P3_Flush    0b0)) ;1729
                                    P1_P1_P3_More = 1'b0; $display(";A 1730");		//(= P1_P1_P3_More    0b0)) ;1730
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 1731");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b11000000)) ;1731
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 1732");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;1732
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 1733");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;1733
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1734");		//(= P1_P1_P3_Flush    0b0)) ;1734
                                    P1_P1_P3_More = 1'b0; $display(";A 1735");		//(= P1_P1_P3_More    0b0)) ;1735
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 1736");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b01000000)) ;1736
                                    P1_P1_P3_EAX <= #1 (P1_P1_P3_EAX + 32'sb00000000000000000000000000000001); $display(";A 1737");		//(= P1_P1_P3_EAX    (bv-add P1_P1_P3_EAX  0b00000000000000000000000000000001))) ;1737
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1738");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1738
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1739");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1739
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1740");		//(= P1_P1_P3_Flush    0b0)) ;1740
                                    P1_P1_P3_More = 1'b0; $display(";A 1741");		//(= P1_P1_P3_More    0b0)) ;1741
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 1742");		//(= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr )   0b01000011)) ;1742
                                    P1_P1_P3_EBX <= #1 (P1_P1_P3_EBX + 32'sb00000000000000000000000000000001); $display(";A 1743");		//(= P1_P1_P3_EBX    (bv-add P1_P1_P3_EBX  0b00000000000000000000000000000001))) ;1743
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1744");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1744
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1745");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1745
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1746");		//(= P1_P1_P3_Flush    0b0)) ;1746
                                    P1_P1_P3_More = 1'b0; $display(";A 1747");		//(= P1_P1_P3_More    0b0)) ;1747
                                end
                            default:
                                begin
                                    $display(";A 1748");		//(= (and (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b10010000) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b01100110) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b11101011) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b11101001) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b11101010) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b10110000) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b10111000) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b10111011) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b10001011) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b10001001) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b11100100) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b11100110) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b00000100) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b00000101) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b11010000) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b11000000) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b01000000) (/= ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ) 0b01000011))   true)) ;1748
                                    P1_P1_P3_InstAddrPointer = (P1_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 1749");		//(= P1_P1_P3_InstAddrPointer    (bv-add P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;1749
                                    P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1750");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1750
                                    P1_P1_P3_Flush = 1'b0; $display(";A 1751");		//(= P1_P1_P3_Flush    0b0)) ;1751
                                    P1_P1_P3_More = 1'b0; $display(";A 1752");		//(= P1_P1_P3_More    0b0)) ;1752
                                end
                        endcase
                        if (((~(P1_P1_P3_InstQueueRd_Addr < P1_P1_P3_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P1_P1_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P1_P1_P3_Flush) | P1_P1_P3_More))) begin
                            $display(";A 1753");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P1_P3_InstQueueRd_Addr  P1_P1_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P1_P3_Flush ) P1_P1_P3_More ))   0b1)) ;1753
                            P1_P1_P3_State2 = 4'sb0111; $display(";A 1755");		//(= P1_P1_P3_State2    0b0111)) ;1755
                        end
                        else begin
                            $display(";A 1754");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P1_P3_InstQueueRd_Addr  P1_P1_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P1_P3_Flush ) P1_P1_P3_More ))   0b0)) ;1754
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 1756");		//(= P1_P1_P3_State2    0b0110)) ;1756
                        P1_P1_P3_Datao <= #1 ((P1_P1_P3_uWord * 32'b00000000000000010000000000000000) + P1_P1_P3_lWord); $display(";A 1757");		//(= P1_P1_P3_Datao    (bv-add (bv-mul P1_P1_P3_uWord  0b00000000000000010000000000000000) P1_P1_P3_lWord ))) ;1757
                        if ((P1_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 1758");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b1)) ;1758
                            P1_P1_P3_RequestPending <= #1 1'b0; $display(";A 1760");		//(= P1_P1_P3_RequestPending    0b0)) ;1760
                            P1_P1_P3_State2 = 4'sb0101; $display(";A 1761");		//(= P1_P1_P3_State2    0b0101)) ;1761
                        end
                        else begin
                            $display(";A 1759");		//(= (bv-comp P1_P1_P3_READY_n  0b0)   0b0)) ;1759
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 1762");		//(= P1_P1_P3_State2    0b0111)) ;1762
                        if (P1_P1_P3_Flush) begin
                            $display(";A 1763");		//(= P1_P1_P3_Flush    0b1)) ;1763
                            P1_P1_P3_InstQueueRd_Addr = 5'sb00001; $display(";A 1765");		//(= P1_P1_P3_InstQueueRd_Addr    0b00001)) ;1765
                            P1_P1_P3_InstQueueWr_Addr = 5'sb00001; $display(";A 1766");		//(= P1_P1_P3_InstQueueWr_Addr    0b00001)) ;1766
                            if ((P1_P1_P3_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 1767");		//(= (bool-to-bv (bv-slt P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;1767
                                P1_P1_P3_fWord = (-P1_P1_P3_InstAddrPointer); $display(";A 1769");		//(= P1_P1_P3_fWord    (bv-neg P1_P1_P3_InstAddrPointer ))) ;1769
                            end
                            else begin
                                $display(";A 1768");		//(= (bool-to-bv (bv-slt P1_P1_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;1768
                                P1_P1_P3_fWord = P1_P1_P3_InstAddrPointer; $display(";A 1770");		//(= P1_P1_P3_fWord    P1_P1_P3_InstAddrPointer )) ;1770
                            end
                            if (((P1_P1_P3_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 1771");		//(= (bv-comp (bv-smod P1_P1_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;1771
                                P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + (P1_P1_P3_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 1773");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  (bv-smod P1_P1_P3_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;1773
                            end
                            else begin
                                $display(";A 1772");		//(= (bv-comp (bv-smod P1_P1_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;1772
                            end
                        end
                        else begin
                            $display(";A 1764");		//(= P1_P1_P3_Flush    0b0)) ;1764
                        end
                        if (((32'b00000000000000000000000000001111 - P1_P1_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 1774");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;1774
                            P1_P1_P3_State2 = 4'sb1000; $display(";A 1776");		//(= P1_P1_P3_State2    0b1000)) ;1776
                            P1_P1_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 1777");		//(= P1_P1_P3_InstQueueWr_Addr    0b00000)) ;1777
                        end
                        else begin
                            $display(";A 1775");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;1775
                            P1_P1_P3_State2 = 4'sb1001; $display(";A 1778");		//(= P1_P1_P3_State2    0b1001)) ;1778
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 1779");		//(= P1_P1_P3_State2    0b1000)) ;1779
                        if ((P1_P1_P3_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 1780");		//(= (bool-to-bv (bv-le P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;1780
                            P1_P1_P3_InstQueue[P1_P1_P3_InstQueueWr_Addr] = P1_P1_P3_InstQueue[P1_P1_P3_InstQueueRd_Addr]; $display(";A 1782");		//(= P1_P1_P3_InstQueue    ( P1_P1_P3_InstQueue P1_P1_P3_InstQueueRd_Addr ))) ;1782
                            P1_P1_P3_InstQueueRd_Addr = ((P1_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1783");		//(= P1_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1783
                            P1_P1_P3_InstQueueWr_Addr = ((P1_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 1784");		//(= P1_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;1784
                            P1_P1_P3_State2 = 4'sb1000; $display(";A 1785");		//(= P1_P1_P3_State2    0b1000)) ;1785
                        end
                        else begin
                            $display(";A 1781");		//(= (bool-to-bv (bv-le P1_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;1781
                            P1_P1_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 1786");		//(= P1_P1_P3_InstQueueRd_Addr    0b00000)) ;1786
                            P1_P1_P3_State2 = 4'sb1001; $display(";A 1787");		//(= P1_P1_P3_State2    0b1001)) ;1787
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 1788");		//(= P1_P1_P3_State2    0b1001)) ;1788
                        P1_P1_P3_rEIP <= #1 P1_P1_P3_PhyAddrPointer; $display(";A 1789");		//(= P1_P1_P3_rEIP    P1_P1_P3_PhyAddrPointer )) ;1789
                        P1_P1_P3_State2 = 4'sb0001; $display(";A 1790");		//(= P1_P1_P3_State2    0b0001)) ;1790
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2469
    always @(posedge P1_P1_P3_RESET or posedge P1_P1_P3_CLOCK) begin
        if ((P1_P1_P3_RESET == 1'b1)) begin
            $display(";A 1791");		//(= (bv-comp P1_P1_P3_RESET  0b1)   0b1)) ;1791
            P1_P1_P3_ByteEnable <= #1 4'b0000; $display(";A 1793");		//(= P1_P1_P3_ByteEnable    0b0000)) ;1793
            P1_P1_P3_NonAligned <= #1 1'b0; $display(";A 1794");		//(= P1_P1_P3_NonAligned    0b0)) ;1794
        end
        else begin
            $display(";A 1792");		//(= (bv-comp P1_P1_P3_RESET  0b1)   0b0)) ;1792
            case (P1_P1_P3_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 1795");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000000)) ;1795
                        case ((P1_P1_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 1796");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;1796
                                    P1_P1_P3_ByteEnable <= #1 4'b1110; $display(";A 1797");		//(= P1_P1_P3_ByteEnable    0b1110)) ;1797
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 1798");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;1798
                                    P1_P1_P3_ByteEnable <= #1 4'b1101; $display(";A 1799");		//(= P1_P1_P3_ByteEnable    0b1101)) ;1799
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 1800");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;1800
                                    P1_P1_P3_ByteEnable <= #1 4'b1011; $display(";A 1801");		//(= P1_P1_P3_ByteEnable    0b1011)) ;1801
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 1802");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;1802
                                    P1_P1_P3_ByteEnable <= #1 4'b0111; $display(";A 1803");		//(= P1_P1_P3_ByteEnable    0b0111)) ;1803
                                end
                            default:
                                begin
                                    $display(";A 1804");		//(= (and (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;1804
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 1805");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000001)) ;1805
                        case ((P1_P1_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 1806");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;1806
                                    P1_P1_P3_ByteEnable <= #1 4'b1100; $display(";A 1807");		//(= P1_P1_P3_ByteEnable    0b1100)) ;1807
                                    P1_P1_P3_NonAligned <= #1 1'b0; $display(";A 1808");		//(= P1_P1_P3_NonAligned    0b0)) ;1808
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 1809");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;1809
                                    P1_P1_P3_ByteEnable <= #1 4'b1001; $display(";A 1810");		//(= P1_P1_P3_ByteEnable    0b1001)) ;1810
                                    P1_P1_P3_NonAligned <= #1 1'b0; $display(";A 1811");		//(= P1_P1_P3_NonAligned    0b0)) ;1811
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 1812");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;1812
                                    P1_P1_P3_ByteEnable <= #1 4'b0011; $display(";A 1813");		//(= P1_P1_P3_ByteEnable    0b0011)) ;1813
                                    P1_P1_P3_NonAligned <= #1 1'b0; $display(";A 1814");		//(= P1_P1_P3_NonAligned    0b0)) ;1814
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 1815");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;1815
                                    P1_P1_P3_ByteEnable <= #1 4'b0111; $display(";A 1816");		//(= P1_P1_P3_ByteEnable    0b0111)) ;1816
                                    P1_P1_P3_NonAligned <= #1 1'b1; $display(";A 1817");		//(= P1_P1_P3_NonAligned    0b1)) ;1817
                                end
                            default:
                                begin
                                    $display(";A 1818");		//(= (and (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;1818
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 1819");		//(= P1_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;1819
                        case ((P1_P1_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 1820");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;1820
                                    P1_P1_P3_ByteEnable <= #1 4'b0000; $display(";A 1821");		//(= P1_P1_P3_ByteEnable    0b0000)) ;1821
                                    P1_P1_P3_NonAligned <= #1 1'b0; $display(";A 1822");		//(= P1_P1_P3_NonAligned    0b0)) ;1822
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 1823");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;1823
                                    P1_P1_P3_ByteEnable <= #1 4'b0001; $display(";A 1824");		//(= P1_P1_P3_ByteEnable    0b0001)) ;1824
                                    P1_P1_P3_NonAligned <= #1 1'b1; $display(";A 1825");		//(= P1_P1_P3_NonAligned    0b1)) ;1825
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 1826");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;1826
                                    P1_P1_P3_NonAligned <= #1 1'b1; $display(";A 1827");		//(= P1_P1_P3_NonAligned    0b1)) ;1827
                                    P1_P1_P3_ByteEnable <= #1 4'b0011; $display(";A 1828");		//(= P1_P1_P3_ByteEnable    0b0011)) ;1828
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 1829");		//(= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;1829
                                    P1_P1_P3_NonAligned <= #1 1'b1; $display(";A 1830");		//(= P1_P1_P3_NonAligned    0b1)) ;1830
                                    P1_P1_P3_ByteEnable <= #1 4'b0111; $display(";A 1831");		//(= P1_P1_P3_ByteEnable    0b0111)) ;1831
                                end
                            default:
                                begin
                                    $display(";A 1832");		//(= (and (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;1832
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 1833");		//(= (and (/= P1_P1_P3_DataWidth  0b00000000000000000000000000000000) (/= P1_P1_P3_DataWidth  0b00000000000000000000000000000001) (/= P1_P1_P3_DataWidth  0b00000000000000000000000000000010))   true)) ;1833
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2615
    always @(posedge P1_P2_reset or posedge P1_P2_clock) begin
        if ((P1_P2_reset == 1'b1)) begin
            P1_P2_buf1 <= #1 32'sb00000000000000000000000000000000; $display(";A 1836");		//(= P1_P2_buf1    0b00000000000000000000000000000000)) ;1836
            P1_P2_ready11 <= #1 1'b0; $display(";A 1837");		//(= P1_P2_ready11    0b0)) ;1837
            P1_P2_ready12 <= #1 1'b0; $display(";A 1838");		//(= P1_P2_ready12    0b0)) ;1838
        end
        else begin
            if (((((((P1_P2_addr1 > 30'b100000000000000000000000000000) & (P1_P2_ads1 == 1'b0)) & (P1_P2_mio1 == 1'b1)) & (P1_P2_dc1 == 1'b0)) & (P1_P2_wr1 == 1'b1)) & (P1_P2_be1 == 4'b0000))) begin
                $display(";A 1839");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P2_addr1  0b100000000000000000000000000000)) (bv-comp P1_P2_ads1  0b0)) (bv-comp P1_P2_mio1  0b1)) (bv-comp P1_P2_dc1  0b0)) (bv-comp P1_P2_wr1  0b1)) (bv-comp P1_P2_be1  0b0000))   0b1)) ;1839
                P1_P2_buf1 <= #1 P1_P2_do1; $display(";A 1841");		//(= P1_P2_buf1    P1_P2_do1 )) ;1841
                P1_P2_ready11 <= #1 1'b0; $display(";A 1842");		//(= P1_P2_ready11    0b0)) ;1842
                P1_P2_ready12 <= #1 1'b1; $display(";A 1843");		//(= P1_P2_ready12    0b1)) ;1843
            end
            else begin
                $display(";A 1840");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P2_addr1  0b100000000000000000000000000000)) (bv-comp P1_P2_ads1  0b0)) (bv-comp P1_P2_mio1  0b1)) (bv-comp P1_P2_dc1  0b0)) (bv-comp P1_P2_wr1  0b1)) (bv-comp P1_P2_be1  0b0000))   0b0)) ;1840
                if (((((((P1_P2_addr2 > 30'b100000000000000000000000000000) & (P1_P2_ads2 == 1'b0)) & (P1_P2_mio2 == 1'b1)) & (P1_P2_dc2 == 1'b0)) & (P1_P2_wr2 == 1'b1)) & (P1_P2_be2 == 4'b0000))) begin
                    $display(";A 1844");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P2_addr2  0b100000000000000000000000000000)) (bv-comp P1_P2_ads2  0b0)) (bv-comp P1_P2_mio2  0b1)) (bv-comp P1_P2_dc2  0b0)) (bv-comp P1_P2_wr2  0b1)) (bv-comp P1_P2_be2  0b0000))   0b1)) ;1844
                    P1_P2_buf1 <= #1 P1_P2_do2; $display(";A 1846");		//(= P1_P2_buf1    P1_P2_do2 )) ;1846
                    P1_P2_ready11 <= #1 1'b1; $display(";A 1847");		//(= P1_P2_ready11    0b1)) ;1847
                    P1_P2_ready12 <= #1 1'b0; $display(";A 1848");		//(= P1_P2_ready12    0b0)) ;1848
                end
                else begin
                    $display(";A 1845");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P1_P2_addr2  0b100000000000000000000000000000)) (bv-comp P1_P2_ads2  0b0)) (bv-comp P1_P2_mio2  0b1)) (bv-comp P1_P2_dc2  0b0)) (bv-comp P1_P2_wr2  0b1)) (bv-comp P1_P2_be2  0b0000))   0b0)) ;1845
                    P1_P2_ready11 <= #1 1'b1; $display(";A 1849");		//(= P1_P2_ready11    0b1)) ;1849
                    P1_P2_ready12 <= #1 1'b1; $display(";A 1850");		//(= P1_P2_ready12    0b1)) ;1850
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2644
    always @(posedge P1_P2_reset or posedge P1_P2_clock) begin
        if ((P1_P2_reset == 1'b1)) begin
            P1_P2_buf2 <= #1 32'sb00000000000000000000000000000000; $display(";A 1853");		//(= P1_P2_buf2    0b00000000000000000000000000000000)) ;1853
            P1_P2_ready21 <= #1 1'b0; $display(";A 1854");		//(= P1_P2_ready21    0b0)) ;1854
            P1_P2_ready22 <= #1 1'b0; $display(";A 1855");		//(= P1_P2_ready22    0b0)) ;1855
        end
        else begin
            if (((((((P1_P2_addr2 < 30'b100000000000000000000000000000) & (P1_P2_ads2 == 1'b0)) & (P1_P2_mio2 == 1'b1)) & (P1_P2_dc2 == 1'b0)) & (P1_P2_wr2 == 1'b1)) & (P1_P2_be2 == 4'b0000))) begin
                $display(";A 1856");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P1_P2_addr2  0b100000000000000000000000000000)) (bv-comp P1_P2_ads2  0b0)) (bv-comp P1_P2_mio2  0b1)) (bv-comp P1_P2_dc2  0b0)) (bv-comp P1_P2_wr2  0b1)) (bv-comp P1_P2_be2  0b0000))   0b1)) ;1856
                P1_P2_buf2 <= #1 P1_P2_do2; $display(";A 1858");		//(= P1_P2_buf2    P1_P2_do2 )) ;1858
                P1_P2_ready21 <= #1 1'b0; $display(";A 1859");		//(= P1_P2_ready21    0b0)) ;1859
                P1_P2_ready22 <= #1 1'b1; $display(";A 1860");		//(= P1_P2_ready22    0b1)) ;1860
            end
            else begin
                $display(";A 1857");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P1_P2_addr2  0b100000000000000000000000000000)) (bv-comp P1_P2_ads2  0b0)) (bv-comp P1_P2_mio2  0b1)) (bv-comp P1_P2_dc2  0b0)) (bv-comp P1_P2_wr2  0b1)) (bv-comp P1_P2_be2  0b0000))   0b0)) ;1857
                if ((((((P1_P2_ads3 == 1'b0) & (P1_P2_mio3 == 1'b1)) & (P1_P2_dc3 == 1'b0)) & (P1_P2_wr3 == 1'b0)) & (P1_P2_be3 == 4'b0000))) begin
                    $display(";A 1861");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P1_P2_ads3  0b0) (bv-comp P1_P2_mio3  0b1)) (bv-comp P1_P2_dc3  0b0)) (bv-comp P1_P2_wr3  0b0)) (bv-comp P1_P2_be3  0b0000))   0b1)) ;1861
                    P1_P2_ready21 <= #1 1'b1; $display(";A 1863");		//(= P1_P2_ready21    0b1)) ;1863
                    P1_P2_ready22 <= #1 1'b0; $display(";A 1864");		//(= P1_P2_ready22    0b0)) ;1864
                end
                else begin
                    $display(";A 1862");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P1_P2_ads3  0b0) (bv-comp P1_P2_mio3  0b1)) (bv-comp P1_P2_dc3  0b0)) (bv-comp P1_P2_wr3  0b0)) (bv-comp P1_P2_be3  0b0000))   0b0)) ;1862
                    P1_P2_ready21 <= #1 1'b1; $display(";A 1865");		//(= P1_P2_ready21    0b1)) ;1865
                    P1_P2_ready22 <= #1 1'b1; $display(";A 1866");		//(= P1_P2_ready22    0b1)) ;1866
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2672
    always @(P1_P2_datai or P1_P2_buf1 or P1_P2_addr1) begin
        if ((P1_P2_addr1 > 30'b100000000000000000000000000000)) begin
            $display(";A 1867");		//(= (bool-to-bv (bv-gt P1_P2_addr1  0b100000000000000000000000000000))   0b1)) ;1867
            P1_P2_di1 <= #1 P1_P2_buf1; $display(";A 1869");		//(= P1_P2_di1    P1_P2_buf1 )) ;1869
        end
        else begin
            $display(";A 1868");		//(= (bool-to-bv (bv-gt P1_P2_addr1  0b100000000000000000000000000000))   0b0)) ;1868
            P1_P2_di1 <= #1 P1_P2_datai; $display(";A 1870");		//(= P1_P2_di1    P1_P2_datai )) ;1870
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2678
    always @(P1_P2_buf2 or P1_P2_buf1 or P1_P2_addr2) begin
        if ((P1_P2_addr2 > 30'b100000000000000000000000000000)) begin
            $display(";A 1871");		//(= (bool-to-bv (bv-gt P1_P2_addr2  0b100000000000000000000000000000))   0b1)) ;1871
            P1_P2_di2 <= #1 P1_P2_buf1; $display(";A 1873");		//(= P1_P2_di2    P1_P2_buf1 )) ;1873
        end
        else begin
            $display(";A 1872");		//(= (bool-to-bv (bv-gt P1_P2_addr2  0b100000000000000000000000000000))   0b0)) ;1872
            P1_P2_di2 <= #1 P1_P2_buf2; $display(";A 1874");		//(= P1_P2_di2    P1_P2_buf2 )) ;1874
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2684
    always @(P1_P2_do3 or P1_P2_do2 or P1_P2_do1 or P1_P2_addr3 or P1_P2_addr2) begin
        if ((((P1_P2_do1 < 32'b00000000000000000000000000000000) & (P1_P2_do2 < 32'b00000000000000000000000000000000)) & (P1_P2_do3 < 32'b00000000000000000000000000000000))) begin
            $display(";A 1875");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P1_P2_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P1_P2_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P1_P2_do3  0b00000000000000000000000000000000)))   0b1)) ;1875
            P1_P2_address2 <= #1 P1_P2_addr3; $display(";A 1877");		//(= P1_P2_address2    P1_P2_addr3 )) ;1877
        end
        else begin
            $display(";A 1876");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P1_P2_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P1_P2_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P1_P2_do3  0b00000000000000000000000000000000)))   0b0)) ;1876
            P1_P2_address2 <= #1 P1_P2_addr2; $display(";A 1878");		//(= P1_P2_address2    P1_P2_addr2 )) ;1878
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2690
    always @(P1_P2_ready22 or P1_P2_ready21 or P1_P2_ready12 or P1_P2_ready11 or P1_P2_ready2 or P1_P2_ready1 or P1_P2_ads3 or P1_P2_ads1 or P1_P2_mio3 or P1_P2_dc3 or P1_P2_wr3 or P1_P2_addr1 or P1_P2_do3 or P1_P2_buf2) begin
        P1_P2_di3 <= #1 P1_P2_buf2; $display(";A 1879");		//(= P1_P2_di3    P1_P2_buf2 )) ;1879
        P1_P2_datao <= #1 P1_P2_do3; $display(";A 1880");		//(= P1_P2_datao    P1_P2_do3 )) ;1880
        P1_P2_address1 <= #1 P1_P2_addr1; $display(";A 1881");		//(= P1_P2_address1    P1_P2_addr1 )) ;1881
        P1_P2_wr <= #1 P1_P2_wr3; $display(";A 1882");		//(= P1_P2_wr    P1_P2_wr3 )) ;1882
        P1_P2_dc <= #1 P1_P2_dc3; $display(";A 1883");		//(= P1_P2_dc    P1_P2_dc3 )) ;1883
        P1_P2_mio <= #1 P1_P2_mio3; $display(";A 1884");		//(= P1_P2_mio    P1_P2_mio3 )) ;1884
        P1_P2_ast1 <= #1 P1_P2_ads1; $display(";A 1885");		//(= P1_P2_ast1    P1_P2_ads1 )) ;1885
        P1_P2_ast2 <= #1 P1_P2_ads3; $display(";A 1886");		//(= P1_P2_ast2    P1_P2_ads3 )) ;1886
        P1_P2_rdy1 <= #1 (P1_P2_ready11 & P1_P2_ready1); $display(";A 1887");		//(= P1_P2_rdy1    (bv-and P1_P2_ready11  P1_P2_ready1 ))) ;1887
        P1_P2_rdy2 <= #1 (P1_P2_ready12 & P1_P2_ready21); $display(";A 1888");		//(= P1_P2_rdy2    (bv-and P1_P2_ready12  P1_P2_ready21 ))) ;1888
        P1_P2_rdy3 <= #1 (P1_P2_ready22 & P1_P2_ready2); $display(";A 1889");		//(= P1_P2_rdy3    (bv-and P1_P2_ready22  P1_P2_ready2 ))) ;1889
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2815
    always @(posedge P1_P2_P1_RESET or posedge P1_P2_P1_CLOCK) begin
        if ((P1_P2_P1_RESET == 1'b1)) begin
            $display(";A 1890");		//(= (bv-comp P1_P2_P1_RESET  0b1)   0b1)) ;1890
            P1_P2_P1_BE_n <= #1 4'b0000; $display(";A 1892");		//(= P1_P2_P1_BE_n    0b0000)) ;1892
            P1_P2_P1_Address <= #1 30'sb000000000000000000000000000000; $display(";A 1893");		//(= P1_P2_P1_Address    0b000000000000000000000000000000)) ;1893
            P1_P2_P1_W_R_n <= #1 1'b0; $display(";A 1894");		//(= P1_P2_P1_W_R_n    0b0)) ;1894
            P1_P2_P1_D_C_n <= #1 1'b0; $display(";A 1895");		//(= P1_P2_P1_D_C_n    0b0)) ;1895
            P1_P2_P1_M_IO_n <= #1 1'b0; $display(";A 1896");		//(= P1_P2_P1_M_IO_n    0b0)) ;1896
            P1_P2_P1_ADS_n <= #1 1'b0; $display(";A 1897");		//(= P1_P2_P1_ADS_n    0b0)) ;1897
            P1_P2_P1_State <= #1 3'sb000; $display(";A 1898");		//(= P1_P2_P1_State    0b000)) ;1898
            P1_P2_P1_StateNA <= #1 1'b0; $display(";A 1899");		//(= P1_P2_P1_StateNA    0b0)) ;1899
            P1_P2_P1_StateBS16 <= #1 1'b0; $display(";A 1900");		//(= P1_P2_P1_StateBS16    0b0)) ;1900
            P1_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 1901");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000000)) ;1901
        end
        else begin
            $display(";A 1891");		//(= (bv-comp P1_P2_P1_RESET  0b1)   0b0)) ;1891
            case (P1_P2_P1_State)
                3'b000 :
                    begin
                        $display(";A 1902");		//(= P1_P2_P1_State    0b000)) ;1902
                        P1_P2_P1_D_C_n <= #1 1'b1; $display(";A 1903");		//(= P1_P2_P1_D_C_n    0b1)) ;1903
                        P1_P2_P1_ADS_n <= #1 1'b1; $display(";A 1904");		//(= P1_P2_P1_ADS_n    0b1)) ;1904
                        P1_P2_P1_State <= #1 3'sb001; $display(";A 1905");		//(= P1_P2_P1_State    0b001)) ;1905
                        P1_P2_P1_StateNA <= #1 1'b1; $display(";A 1906");		//(= P1_P2_P1_StateNA    0b1)) ;1906
                        P1_P2_P1_StateBS16 <= #1 1'b1; $display(";A 1907");		//(= P1_P2_P1_StateBS16    0b1)) ;1907
                        P1_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 1908");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;1908
                        P1_P2_P1_State <= #1 3'sb001; $display(";A 1909");		//(= P1_P2_P1_State    0b001)) ;1909
                    end
                3'b001 :
                    begin
                        $display(";A 1910");		//(= P1_P2_P1_State    0b001)) ;1910
                        if ((P1_P2_P1_RequestPending == 1'b1)) begin
                            $display(";A 1911");		//(= (bv-comp P1_P2_P1_RequestPending  0b1)   0b1)) ;1911
                            P1_P2_P1_State <= #1 3'sb010; $display(";A 1913");		//(= P1_P2_P1_State    0b010)) ;1913
                        end
                        else begin
                            $display(";A 1912");		//(= (bv-comp P1_P2_P1_RequestPending  0b1)   0b0)) ;1912
                            if ((P1_P2_P1_HOLD == 1'b1)) begin
                                $display(";A 1914");		//(= (bv-comp P1_P2_P1_HOLD  0b1)   0b1)) ;1914
                                P1_P2_P1_State <= #1 3'sb101; $display(";A 1916");		//(= P1_P2_P1_State    0b101)) ;1916
                            end
                            else begin
                                $display(";A 1915");		//(= (bv-comp P1_P2_P1_HOLD  0b1)   0b0)) ;1915
                                P1_P2_P1_State <= #1 3'sb001; $display(";A 1917");		//(= P1_P2_P1_State    0b001)) ;1917
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 1918");		//(= P1_P2_P1_State    0b010)) ;1918
                        P1_P2_P1_Address <= #1 ((P1_P2_P1_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 1919");		//(= P1_P2_P1_Address    (bv-smod (bv-sdiv P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;1919
                        P1_P2_P1_BE_n <= #1 P1_P2_P1_ByteEnable; $display(";A 1920");		//(= P1_P2_P1_BE_n    P1_P2_P1_ByteEnable )) ;1920
                        P1_P2_P1_M_IO_n <= #1 P1_P2_P1_MemoryFetch; $display(";A 1921");		//(= P1_P2_P1_M_IO_n    P1_P2_P1_MemoryFetch )) ;1921
                        if ((P1_P2_P1_ReadRequest == 1'b1)) begin
                            $display(";A 1922");		//(= (bv-comp P1_P2_P1_ReadRequest  0b1)   0b1)) ;1922
                            P1_P2_P1_W_R_n <= #1 1'b0; $display(";A 1924");		//(= P1_P2_P1_W_R_n    0b0)) ;1924
                        end
                        else begin
                            $display(";A 1923");		//(= (bv-comp P1_P2_P1_ReadRequest  0b1)   0b0)) ;1923
                            P1_P2_P1_W_R_n <= #1 1'b1; $display(";A 1925");		//(= P1_P2_P1_W_R_n    0b1)) ;1925
                        end
                        if ((P1_P2_P1_CodeFetch == 1'b1)) begin
                            $display(";A 1926");		//(= (bv-comp P1_P2_P1_CodeFetch  0b1)   0b1)) ;1926
                            P1_P2_P1_D_C_n <= #1 1'b0; $display(";A 1928");		//(= P1_P2_P1_D_C_n    0b0)) ;1928
                        end
                        else begin
                            $display(";A 1927");		//(= (bv-comp P1_P2_P1_CodeFetch  0b1)   0b0)) ;1927
                            P1_P2_P1_D_C_n <= #1 1'b1; $display(";A 1929");		//(= P1_P2_P1_D_C_n    0b1)) ;1929
                        end
                        P1_P2_P1_ADS_n <= #1 1'b0; $display(";A 1930");		//(= P1_P2_P1_ADS_n    0b0)) ;1930
                        P1_P2_P1_State <= #1 3'sb011; $display(";A 1931");		//(= P1_P2_P1_State    0b011)) ;1931
                    end
                3'b011 :
                    begin
                        $display(";A 1932");		//(= P1_P2_P1_State    0b011)) ;1932
                        if ((((P1_P2_P1_READY_n == 1'b0) & (P1_P2_P1_HOLD == 1'b0)) & (P1_P2_P1_RequestPending == 1'b1))) begin
                            $display(";A 1933");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b1))   0b1)) ;1933
                            P1_P2_P1_State <= #1 3'sb010; $display(";A 1935");		//(= P1_P2_P1_State    0b010)) ;1935
                        end
                        else begin
                            $display(";A 1934");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b1))   0b0)) ;1934
                            if (((P1_P2_P1_READY_n == 1'b1) & (P1_P2_P1_NA_n == 1'b1))) begin
                                $display(";A 1936");		//(= (bv-and (bv-comp P1_P2_P1_READY_n  0b1) (bv-comp P1_P2_P1_NA_n  0b1))   0b1)) ;1936
                            end
                            else begin
                                $display(";A 1937");		//(= (bv-and (bv-comp P1_P2_P1_READY_n  0b1) (bv-comp P1_P2_P1_NA_n  0b1))   0b0)) ;1937
                                if ((((P1_P2_P1_RequestPending == 1'b1) | (P1_P2_P1_HOLD == 1'b1)) & ((P1_P2_P1_READY_n == 1'b1) & (P1_P2_P1_NA_n == 1'b0)))) begin
                                    $display(";A 1938");		//(= (bv-and (bv-or (bv-comp P1_P2_P1_RequestPending  0b1) (bv-comp P1_P2_P1_HOLD  0b1)) (bv-and (bv-comp P1_P2_P1_READY_n  0b1) (bv-comp P1_P2_P1_NA_n  0b0)))   0b1)) ;1938
                                    P1_P2_P1_State <= #1 3'sb111; $display(";A 1940");		//(= P1_P2_P1_State    0b111)) ;1940
                                end
                                else begin
                                    $display(";A 1939");		//(= (bv-and (bv-or (bv-comp P1_P2_P1_RequestPending  0b1) (bv-comp P1_P2_P1_HOLD  0b1)) (bv-and (bv-comp P1_P2_P1_READY_n  0b1) (bv-comp P1_P2_P1_NA_n  0b0)))   0b0)) ;1939
                                    if (((((P1_P2_P1_RequestPending == 1'b1) & (P1_P2_P1_HOLD == 1'b0)) & (P1_P2_P1_READY_n == 1'b1)) & (P1_P2_P1_NA_n == 1'b0))) begin
                                        $display(";A 1941");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P2_P1_RequestPending  0b1) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_READY_n  0b1)) (bv-comp P1_P2_P1_NA_n  0b0))   0b1)) ;1941
                                        P1_P2_P1_State <= #1 3'sb110; $display(";A 1943");		//(= P1_P2_P1_State    0b110)) ;1943
                                    end
                                    else begin
                                        $display(";A 1942");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P2_P1_RequestPending  0b1) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_READY_n  0b1)) (bv-comp P1_P2_P1_NA_n  0b0))   0b0)) ;1942
                                        if ((((P1_P2_P1_RequestPending == 1'b0) & (P1_P2_P1_HOLD == 1'b0)) & (P1_P2_P1_READY_n == 1'b0))) begin
                                            $display(";A 1944");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_RequestPending  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_READY_n  0b0))   0b1)) ;1944
                                            P1_P2_P1_State <= #1 3'sb001; $display(";A 1946");		//(= P1_P2_P1_State    0b001)) ;1946
                                        end
                                        else begin
                                            $display(";A 1945");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_RequestPending  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_READY_n  0b0))   0b0)) ;1945
                                            if (((P1_P2_P1_HOLD == 1'b1) & (P1_P2_P1_READY_n == 1'b1))) begin
                                                $display(";A 1947");		//(= (bv-and (bv-comp P1_P2_P1_HOLD  0b1) (bv-comp P1_P2_P1_READY_n  0b1))   0b1)) ;1947
                                                P1_P2_P1_State <= #1 3'sb101; $display(";A 1949");		//(= P1_P2_P1_State    0b101)) ;1949
                                            end
                                            else begin
                                                $display(";A 1948");		//(= (bv-and (bv-comp P1_P2_P1_HOLD  0b1) (bv-comp P1_P2_P1_READY_n  0b1))   0b0)) ;1948
                                                P1_P2_P1_State <= #1 3'sb011; $display(";A 1950");		//(= P1_P2_P1_State    0b011)) ;1950
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P1_P2_P1_StateBS16 <= #1 P1_P2_P1_BS16_n; $display(";A 1951");		//(= P1_P2_P1_StateBS16    P1_P2_P1_BS16_n )) ;1951
                        if ((P1_P2_P1_BS16_n == 1'b0)) begin
                            $display(";A 1952");		//(= (bv-comp P1_P2_P1_BS16_n  0b0)   0b1)) ;1952
                            P1_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 1954");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000001)) ;1954
                        end
                        else begin
                            $display(";A 1953");		//(= (bv-comp P1_P2_P1_BS16_n  0b0)   0b0)) ;1953
                            P1_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 1955");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;1955
                        end
                        P1_P2_P1_StateNA <= #1 P1_P2_P1_NA_n; $display(";A 1956");		//(= P1_P2_P1_StateNA    P1_P2_P1_NA_n )) ;1956
                        P1_P2_P1_ADS_n <= #1 1'b1; $display(";A 1957");		//(= P1_P2_P1_ADS_n    0b1)) ;1957
                    end
                3'b100 :
                    begin
                        $display(";A 1958");		//(= P1_P2_P1_State    0b100)) ;1958
                        if ((((P1_P2_P1_NA_n == 1'b0) & (P1_P2_P1_HOLD == 1'b0)) & (P1_P2_P1_RequestPending == 1'b1))) begin
                            $display(";A 1959");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_NA_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b1))   0b1)) ;1959
                            P1_P2_P1_State <= #1 3'sb110; $display(";A 1961");		//(= P1_P2_P1_State    0b110)) ;1961
                        end
                        else begin
                            $display(";A 1960");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_NA_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b1))   0b0)) ;1960
                            if (((P1_P2_P1_NA_n == 1'b0) & ((P1_P2_P1_HOLD == 1'b1) | (P1_P2_P1_RequestPending == 1'b0)))) begin
                                $display(";A 1962");		//(= (bv-and (bv-comp P1_P2_P1_NA_n  0b0) (bv-or (bv-comp P1_P2_P1_HOLD  0b1) (bv-comp P1_P2_P1_RequestPending  0b0)))   0b1)) ;1962
                                P1_P2_P1_State <= #1 3'sb111; $display(";A 1964");		//(= P1_P2_P1_State    0b111)) ;1964
                            end
                            else begin
                                $display(";A 1963");		//(= (bv-and (bv-comp P1_P2_P1_NA_n  0b0) (bv-or (bv-comp P1_P2_P1_HOLD  0b1) (bv-comp P1_P2_P1_RequestPending  0b0)))   0b0)) ;1963
                                if ((P1_P2_P1_NA_n == 1'b1)) begin
                                    $display(";A 1965");		//(= (bv-comp P1_P2_P1_NA_n  0b1)   0b1)) ;1965
                                    P1_P2_P1_State <= #1 3'sb011; $display(";A 1967");		//(= P1_P2_P1_State    0b011)) ;1967
                                end
                                else begin
                                    $display(";A 1966");		//(= (bv-comp P1_P2_P1_NA_n  0b1)   0b0)) ;1966
                                    P1_P2_P1_State <= #1 3'sb100; $display(";A 1968");		//(= P1_P2_P1_State    0b100)) ;1968
                                end
                            end
                        end
                        P1_P2_P1_StateBS16 <= #1 P1_P2_P1_BS16_n; $display(";A 1969");		//(= P1_P2_P1_StateBS16    P1_P2_P1_BS16_n )) ;1969
                        if ((P1_P2_P1_BS16_n == 1'b0)) begin
                            $display(";A 1970");		//(= (bv-comp P1_P2_P1_BS16_n  0b0)   0b1)) ;1970
                            P1_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 1972");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000001)) ;1972
                        end
                        else begin
                            $display(";A 1971");		//(= (bv-comp P1_P2_P1_BS16_n  0b0)   0b0)) ;1971
                            P1_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 1973");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;1973
                        end
                        P1_P2_P1_StateNA <= #1 P1_P2_P1_NA_n; $display(";A 1974");		//(= P1_P2_P1_StateNA    P1_P2_P1_NA_n )) ;1974
                        P1_P2_P1_ADS_n <= #1 1'b1; $display(";A 1975");		//(= P1_P2_P1_ADS_n    0b1)) ;1975
                    end
                3'b101 :
                    begin
                        $display(";A 1976");		//(= P1_P2_P1_State    0b101)) ;1976
                        if (((P1_P2_P1_HOLD == 1'b0) & (P1_P2_P1_RequestPending == 1'b1))) begin
                            $display(";A 1977");		//(= (bv-and (bv-comp P1_P2_P1_HOLD  0b0) (bv-comp P1_P2_P1_RequestPending  0b1))   0b1)) ;1977
                            P1_P2_P1_State <= #1 3'sb010; $display(";A 1979");		//(= P1_P2_P1_State    0b010)) ;1979
                        end
                        else begin
                            $display(";A 1978");		//(= (bv-and (bv-comp P1_P2_P1_HOLD  0b0) (bv-comp P1_P2_P1_RequestPending  0b1))   0b0)) ;1978
                            if (((P1_P2_P1_HOLD == 1'b0) & (P1_P2_P1_RequestPending == 1'b0))) begin
                                $display(";A 1980");		//(= (bv-and (bv-comp P1_P2_P1_HOLD  0b0) (bv-comp P1_P2_P1_RequestPending  0b0))   0b1)) ;1980
                                P1_P2_P1_State <= #1 3'sb001; $display(";A 1982");		//(= P1_P2_P1_State    0b001)) ;1982
                            end
                            else begin
                                $display(";A 1981");		//(= (bv-and (bv-comp P1_P2_P1_HOLD  0b0) (bv-comp P1_P2_P1_RequestPending  0b0))   0b0)) ;1981
                                P1_P2_P1_State <= #1 3'sb101; $display(";A 1983");		//(= P1_P2_P1_State    0b101)) ;1983
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 1984");		//(= P1_P2_P1_State    0b110)) ;1984
                        P1_P2_P1_Address <= #1 ((P1_P2_P1_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 1985");		//(= P1_P2_P1_Address    (bv-smod (bv-sdiv P1_P2_P1_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;1985
                        P1_P2_P1_BE_n <= #1 P1_P2_P1_ByteEnable; $display(";A 1986");		//(= P1_P2_P1_BE_n    P1_P2_P1_ByteEnable )) ;1986
                        P1_P2_P1_M_IO_n <= #1 P1_P2_P1_MemoryFetch; $display(";A 1987");		//(= P1_P2_P1_M_IO_n    P1_P2_P1_MemoryFetch )) ;1987
                        if ((P1_P2_P1_ReadRequest == 1'b1)) begin
                            $display(";A 1988");		//(= (bv-comp P1_P2_P1_ReadRequest  0b1)   0b1)) ;1988
                            P1_P2_P1_W_R_n <= #1 1'b0; $display(";A 1990");		//(= P1_P2_P1_W_R_n    0b0)) ;1990
                        end
                        else begin
                            $display(";A 1989");		//(= (bv-comp P1_P2_P1_ReadRequest  0b1)   0b0)) ;1989
                            P1_P2_P1_W_R_n <= #1 1'b1; $display(";A 1991");		//(= P1_P2_P1_W_R_n    0b1)) ;1991
                        end
                        if ((P1_P2_P1_CodeFetch == 1'b1)) begin
                            $display(";A 1992");		//(= (bv-comp P1_P2_P1_CodeFetch  0b1)   0b1)) ;1992
                            P1_P2_P1_D_C_n <= #1 1'b0; $display(";A 1994");		//(= P1_P2_P1_D_C_n    0b0)) ;1994
                        end
                        else begin
                            $display(";A 1993");		//(= (bv-comp P1_P2_P1_CodeFetch  0b1)   0b0)) ;1993
                            P1_P2_P1_D_C_n <= #1 1'b1; $display(";A 1995");		//(= P1_P2_P1_D_C_n    0b1)) ;1995
                        end
                        P1_P2_P1_ADS_n <= #1 1'b0; $display(";A 1996");		//(= P1_P2_P1_ADS_n    0b0)) ;1996
                        if ((P1_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 1997");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;1997
                            P1_P2_P1_State <= #1 3'sb100; $display(";A 1999");		//(= P1_P2_P1_State    0b100)) ;1999
                        end
                        else begin
                            $display(";A 1998");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;1998
                            P1_P2_P1_State <= #1 3'sb110; $display(";A 2000");		//(= P1_P2_P1_State    0b110)) ;2000
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 2001");		//(= P1_P2_P1_State    0b111)) ;2001
                        if ((((P1_P2_P1_READY_n == 1'b1) & (P1_P2_P1_RequestPending == 1'b1)) & (P1_P2_P1_HOLD == 1'b0))) begin
                            $display(";A 2002");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b1) (bv-comp P1_P2_P1_RequestPending  0b1)) (bv-comp P1_P2_P1_HOLD  0b0))   0b1)) ;2002
                            P1_P2_P1_State <= #1 3'sb110; $display(";A 2004");		//(= P1_P2_P1_State    0b110)) ;2004
                        end
                        else begin
                            $display(";A 2003");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b1) (bv-comp P1_P2_P1_RequestPending  0b1)) (bv-comp P1_P2_P1_HOLD  0b0))   0b0)) ;2003
                            if (((P1_P2_P1_READY_n == 1'b0) & (P1_P2_P1_HOLD == 1'b1))) begin
                                $display(";A 2005");		//(= (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b1))   0b1)) ;2005
                                P1_P2_P1_State <= #1 3'sb101; $display(";A 2007");		//(= P1_P2_P1_State    0b101)) ;2007
                            end
                            else begin
                                $display(";A 2006");		//(= (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b1))   0b0)) ;2006
                                if ((((P1_P2_P1_READY_n == 1'b0) & (P1_P2_P1_HOLD == 1'b0)) & (P1_P2_P1_RequestPending == 1'b1))) begin
                                    $display(";A 2008");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b1))   0b1)) ;2008
                                    P1_P2_P1_State <= #1 3'sb010; $display(";A 2010");		//(= P1_P2_P1_State    0b010)) ;2010
                                end
                                else begin
                                    $display(";A 2009");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b1))   0b0)) ;2009
                                    if ((((P1_P2_P1_READY_n == 1'b0) & (P1_P2_P1_HOLD == 1'b0)) & (P1_P2_P1_RequestPending == 1'b0))) begin
                                        $display(";A 2011");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b0))   0b1)) ;2011
                                        P1_P2_P1_State <= #1 3'sb001; $display(";A 2013");		//(= P1_P2_P1_State    0b001)) ;2013
                                    end
                                    else begin
                                        $display(";A 2012");		//(= (bv-and (bv-and (bv-comp P1_P2_P1_READY_n  0b0) (bv-comp P1_P2_P1_HOLD  0b0)) (bv-comp P1_P2_P1_RequestPending  0b0))   0b0)) ;2012
                                        P1_P2_P1_State <= #1 3'sb111; $display(";A 2014");		//(= P1_P2_P1_State    0b111)) ;2014
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:2959
    always @(posedge P1_P2_P1_RESET or posedge P1_P2_P1_CLOCK) begin
        if ((P1_P2_P1_RESET == 1'b1)) begin
            $display(";A 2015");		//(= (bv-comp P1_P2_P1_RESET  0b1)   0b1)) ;2015
            P1_P2_P1_State2 = 4'sb0000; $display(";A 2017");		//(= P1_P2_P1_State2    0b0000)) ;2017
            P1_P2_P1_InstQueue[0] = 8'b00000000; $display(";A 2018");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2018
            P1_P2_P1_InstQueue[1] = 8'b00000000; $display(";A 2019");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2019
            P1_P2_P1_InstQueue[2] = 8'b00000000; $display(";A 2020");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2020
            P1_P2_P1_InstQueue[3] = 8'b00000000; $display(";A 2021");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2021
            P1_P2_P1_InstQueue[4] = 8'b00000000; $display(";A 2022");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2022
            P1_P2_P1_InstQueue[5] = 8'b00000000; $display(";A 2023");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2023
            P1_P2_P1_InstQueue[6] = 8'b00000000; $display(";A 2024");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2024
            P1_P2_P1_InstQueue[7] = 8'b00000000; $display(";A 2025");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2025
            P1_P2_P1_InstQueue[8] = 8'b00000000; $display(";A 2026");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2026
            P1_P2_P1_InstQueue[9] = 8'b00000000; $display(";A 2027");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2027
            P1_P2_P1_InstQueue[10] = 8'b00000000; $display(";A 2028");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2028
            P1_P2_P1_InstQueue[11] = 8'b00000000; $display(";A 2029");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2029
            P1_P2_P1_InstQueue[12] = 8'b00000000; $display(";A 2030");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2030
            P1_P2_P1_InstQueue[13] = 8'b00000000; $display(";A 2031");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2031
            P1_P2_P1_InstQueue[14] = 8'b00000000; $display(";A 2032");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2032
            P1_P2_P1_InstQueue[15] = 8'b00000000; $display(";A 2033");		//(= P1_P2_P1_InstQueue    0b00000000)) ;2033
            P1_P2_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 2034");		//(= P1_P2_P1_InstQueueRd_Addr    0b00000)) ;2034
            P1_P2_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 2035");		//(= P1_P2_P1_InstQueueWr_Addr    0b00000)) ;2035
            P1_P2_P1_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 2036");		//(= P1_P2_P1_InstAddrPointer    0b00000000000000000000000000000000)) ;2036
            P1_P2_P1_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 2037");		//(= P1_P2_P1_PhyAddrPointer    0b00000000000000000000000000000000)) ;2037
            P1_P2_P1_Extended = 1'b0; $display(";A 2038");		//(= P1_P2_P1_Extended    0b0)) ;2038
            P1_P2_P1_More = 1'b0; $display(";A 2039");		//(= P1_P2_P1_More    0b0)) ;2039
            P1_P2_P1_Flush = 1'b0; $display(";A 2040");		//(= P1_P2_P1_Flush    0b0)) ;2040
            P1_P2_P1_lWord = 16'sb0000000000000000; $display(";A 2041");		//(= P1_P2_P1_lWord    0b0000000000000000)) ;2041
            P1_P2_P1_uWord = 15'sb000000000000000; $display(";A 2042");		//(= P1_P2_P1_uWord    0b000000000000000)) ;2042
            P1_P2_P1_fWord = 32'sb00000000000000000000000000000000; $display(";A 2043");		//(= P1_P2_P1_fWord    0b00000000000000000000000000000000)) ;2043
            P1_P2_P1_CodeFetch <= #1 1'b0; $display(";A 2044");		//(= P1_P2_P1_CodeFetch    0b0)) ;2044
            P1_P2_P1_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 2045");		//(= P1_P2_P1_Datao    0b00000000000000000000000000000000)) ;2045
            P1_P2_P1_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 2046");		//(= P1_P2_P1_EAX    0b00000000000000000000000000000000)) ;2046
            P1_P2_P1_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 2047");		//(= P1_P2_P1_EBX    0b00000000000000000000000000000000)) ;2047
            P1_P2_P1_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 2048");		//(= P1_P2_P1_rEIP    0b00000000000000000000000000000000)) ;2048
            P1_P2_P1_ReadRequest <= #1 1'b0; $display(";A 2049");		//(= P1_P2_P1_ReadRequest    0b0)) ;2049
            P1_P2_P1_MemoryFetch <= #1 1'b0; $display(";A 2050");		//(= P1_P2_P1_MemoryFetch    0b0)) ;2050
            P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2051");		//(= P1_P2_P1_RequestPending    0b0)) ;2051
        end
        else begin
            $display(";A 2016");		//(= (bv-comp P1_P2_P1_RESET  0b1)   0b0)) ;2016
            case (P1_P2_P1_State2)
                4'b0000 :
                    begin
                        $display(";A 2052");		//(= P1_P2_P1_State2    0b0000)) ;2052
                        P1_P2_P1_PhyAddrPointer = P1_P2_P1_rEIP; $display(";A 2053");		//(= P1_P2_P1_PhyAddrPointer    P1_P2_P1_rEIP )) ;2053
                        P1_P2_P1_InstAddrPointer = P1_P2_P1_PhyAddrPointer; $display(";A 2054");		//(= P1_P2_P1_InstAddrPointer    P1_P2_P1_PhyAddrPointer )) ;2054
                        P1_P2_P1_State2 = 4'sb0001; $display(";A 2055");		//(= P1_P2_P1_State2    0b0001)) ;2055
                        P1_P2_P1_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 2056");		//(= P1_P2_P1_rEIP    0b00000000000011111111111111110000)) ;2056
                        P1_P2_P1_ReadRequest <= #1 1'b1; $display(";A 2057");		//(= P1_P2_P1_ReadRequest    0b1)) ;2057
                        P1_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 2058");		//(= P1_P2_P1_MemoryFetch    0b1)) ;2058
                        P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2059");		//(= P1_P2_P1_RequestPending    0b1)) ;2059
                    end
                4'b0001 :
                    begin
                        $display(";A 2060");		//(= P1_P2_P1_State2    0b0001)) ;2060
                        P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2061");		//(= P1_P2_P1_RequestPending    0b1)) ;2061
                        P1_P2_P1_ReadRequest <= #1 1'b1; $display(";A 2062");		//(= P1_P2_P1_ReadRequest    0b1)) ;2062
                        P1_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 2063");		//(= P1_P2_P1_MemoryFetch    0b1)) ;2063
                        P1_P2_P1_CodeFetch <= #1 1'b1; $display(";A 2064");		//(= P1_P2_P1_CodeFetch    0b1)) ;2064
                        if ((P1_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 2065");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2065
                            P1_P2_P1_State2 = 4'sb0010; $display(";A 2067");		//(= P1_P2_P1_State2    0b0010)) ;2067
                        end
                        else begin
                            $display(";A 2066");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2066
                            P1_P2_P1_State2 = 4'sb0001; $display(";A 2068");		//(= P1_P2_P1_State2    0b0001)) ;2068
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 2069");		//(= P1_P2_P1_State2    0b0010)) ;2069
                        P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2070");		//(= P1_P2_P1_RequestPending    0b0)) ;2070
                        P1_P2_P1_InstQueue[P1_P2_P1_InstQueueWr_Addr] = (P1_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 2071");		//(= P1_P2_P1_InstQueue    (bv-smod P1_P2_P1_Datai  0b00000000000000000000000100000000))) ;2071
                        P1_P2_P1_InstQueueWr_Addr = ((P1_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2072");		//(= P1_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2072
                        P1_P2_P1_InstQueue[P1_P2_P1_InstQueueWr_Addr] = (P1_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 2073");		//(= P1_P2_P1_InstQueue    (bv-smod P1_P2_P1_Datai  0b00000000000000000000000100000000))) ;2073
                        P1_P2_P1_InstQueueWr_Addr = ((P1_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2074");		//(= P1_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2074
                        if ((P1_P2_P1_StateBS16 == 1'b1)) begin
                            $display(";A 2075");		//(= (bv-comp P1_P2_P1_StateBS16  0b1)   0b1)) ;2075
                            P1_P2_P1_InstQueue[P1_P2_P1_InstQueueWr_Addr] = ((P1_P2_P1_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 2077");		//(= P1_P2_P1_InstQueue    (bv-smod (bv-sdiv P1_P2_P1_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;2077
                            P1_P2_P1_InstQueueWr_Addr = ((P1_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2078");		//(= P1_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2078
                            P1_P2_P1_InstQueue[P1_P2_P1_InstQueueWr_Addr] = ((P1_P2_P1_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 2079");		//(= P1_P2_P1_InstQueue    (bv-smod (bv-sdiv P1_P2_P1_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;2079
                            P1_P2_P1_InstQueueWr_Addr = ((P1_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2080");		//(= P1_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2080
                            P1_P2_P1_PhyAddrPointer = (P1_P2_P1_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 2081");		//(= P1_P2_P1_PhyAddrPointer    (bv-add P1_P2_P1_PhyAddrPointer  0b00000000000000000000000000000100))) ;2081
                            P1_P2_P1_State2 = 4'sb0101; $display(";A 2082");		//(= P1_P2_P1_State2    0b0101)) ;2082
                        end
                        else begin
                            $display(";A 2076");		//(= (bv-comp P1_P2_P1_StateBS16  0b1)   0b0)) ;2076
                            P1_P2_P1_PhyAddrPointer = (P1_P2_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2083");		//(= P1_P2_P1_PhyAddrPointer    (bv-add P1_P2_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;2083
                            if ((P1_P2_P1_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 2084");		//(= (bool-to-bv (bv-slt P1_P2_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;2084
                                P1_P2_P1_rEIP <= #1 (-P1_P2_P1_PhyAddrPointer); $display(";A 2086");		//(= P1_P2_P1_rEIP    (bv-neg P1_P2_P1_PhyAddrPointer ))) ;2086
                            end
                            else begin
                                $display(";A 2085");		//(= (bool-to-bv (bv-slt P1_P2_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;2085
                                P1_P2_P1_rEIP <= #1 P1_P2_P1_PhyAddrPointer; $display(";A 2087");		//(= P1_P2_P1_rEIP    P1_P2_P1_PhyAddrPointer )) ;2087
                            end
                            P1_P2_P1_State2 = 4'sb0011; $display(";A 2088");		//(= P1_P2_P1_State2    0b0011)) ;2088
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 2089");		//(= P1_P2_P1_State2    0b0011)) ;2089
                        P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2090");		//(= P1_P2_P1_RequestPending    0b1)) ;2090
                        if ((P1_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 2091");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2091
                            P1_P2_P1_State2 = 4'sb0100; $display(";A 2093");		//(= P1_P2_P1_State2    0b0100)) ;2093
                        end
                        else begin
                            $display(";A 2092");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2092
                            P1_P2_P1_State2 = 4'sb0011; $display(";A 2094");		//(= P1_P2_P1_State2    0b0011)) ;2094
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 2095");		//(= P1_P2_P1_State2    0b0100)) ;2095
                        P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2096");		//(= P1_P2_P1_RequestPending    0b0)) ;2096
                        P1_P2_P1_InstQueue[P1_P2_P1_InstQueueWr_Addr] = (P1_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 2097");		//(= P1_P2_P1_InstQueue    (bv-smod P1_P2_P1_Datai  0b00000000000000000000000100000000))) ;2097
                        P1_P2_P1_InstQueueWr_Addr = ((P1_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2098");		//(= P1_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2098
                        P1_P2_P1_InstQueue[P1_P2_P1_InstQueueWr_Addr] = (P1_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 2099");		//(= P1_P2_P1_InstQueue    (bv-smod P1_P2_P1_Datai  0b00000000000000000000000100000000))) ;2099
                        P1_P2_P1_InstQueueWr_Addr = ((P1_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2100");		//(= P1_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2100
                        P1_P2_P1_PhyAddrPointer = (P1_P2_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2101");		//(= P1_P2_P1_PhyAddrPointer    (bv-add P1_P2_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;2101
                        P1_P2_P1_State2 = 4'sb0101; $display(";A 2102");		//(= P1_P2_P1_State2    0b0101)) ;2102
                    end
                4'b0101 :
                    begin
                        $display(";A 2103");		//(= P1_P2_P1_State2    0b0101)) ;2103
                        case (P1_P2_P1_InstQueue[P1_P2_P1_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 2104");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b10010000)) ;2104
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2105");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2105
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2106");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2106
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2107");		//(= P1_P2_P1_Flush    0b0)) ;2107
                                    P1_P2_P1_More = 1'b0; $display(";A 2108");		//(= P1_P2_P1_More    0b0)) ;2108
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 2109");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b01100110)) ;2109
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2110");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2110
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2111");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2111
                                    P1_P2_P1_Extended = 1'b1; $display(";A 2112");		//(= P1_P2_P1_Extended    0b1)) ;2112
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2113");		//(= P1_P2_P1_Flush    0b0)) ;2113
                                    P1_P2_P1_More = 1'b0; $display(";A 2114");		//(= P1_P2_P1_More    0b0)) ;2114
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 2115");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b11101011)) ;2115
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 2116");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;2116
                                        if ((P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 2118");		//(= (bool-to-bv (bv-gt P1_P2_P1_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;2118
                                            P1_P2_P1_PhyAddrPointer = ((P1_P2_P1_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 2120");		//(= P1_P2_P1_PhyAddrPointer    (bv-sub (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P1_P2_P1_InstQueue 0 )))) ;2120
                                            P1_P2_P1_InstAddrPointer = P1_P2_P1_PhyAddrPointer; $display(";A 2121");		//(= P1_P2_P1_InstAddrPointer    P1_P2_P1_PhyAddrPointer )) ;2121
                                        end
                                        else begin
                                            $display(";A 2119");		//(= (bool-to-bv (bv-gt P1_P2_P1_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;2119
                                            P1_P2_P1_PhyAddrPointer = ((P1_P2_P1_InstAddrPointer + 32'b00000000000000000000000000000010) + P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 2122");		//(= P1_P2_P1_PhyAddrPointer    (bv-add (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000010) P1_P2_P1_InstQueue 0 ))) ;2122
                                            P1_P2_P1_InstAddrPointer = P1_P2_P1_PhyAddrPointer; $display(";A 2123");		//(= P1_P2_P1_InstAddrPointer    P1_P2_P1_PhyAddrPointer )) ;2123
                                        end
                                        P1_P2_P1_Flush = 1'b1; $display(";A 2124");		//(= P1_P2_P1_Flush    0b1)) ;2124
                                        P1_P2_P1_More = 1'b0; $display(";A 2125");		//(= P1_P2_P1_More    0b0)) ;2125
                                    end
                                    else begin
                                        $display(";A 2117");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;2117
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2126");		//(= P1_P2_P1_Flush    0b0)) ;2126
                                        P1_P2_P1_More = 1'b1; $display(";A 2127");		//(= P1_P2_P1_More    0b1)) ;2127
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 2128");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b11101001)) ;2128
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 2129");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;2129
                                        P1_P2_P1_PhyAddrPointer = ((P1_P2_P1_InstAddrPointer + 32'b00000000000000000000000000000101) + P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 2131");		//(= P1_P2_P1_PhyAddrPointer    (bv-add (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000101) P1_P2_P1_InstQueue 0 ))) ;2131
                                        P1_P2_P1_InstAddrPointer = P1_P2_P1_PhyAddrPointer; $display(";A 2132");		//(= P1_P2_P1_InstAddrPointer    P1_P2_P1_PhyAddrPointer )) ;2132
                                        P1_P2_P1_Flush = 1'b1; $display(";A 2133");		//(= P1_P2_P1_Flush    0b1)) ;2133
                                        P1_P2_P1_More = 1'b0; $display(";A 2134");		//(= P1_P2_P1_More    0b0)) ;2134
                                    end
                                    else begin
                                        $display(";A 2130");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;2130
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2135");		//(= P1_P2_P1_Flush    0b0)) ;2135
                                        P1_P2_P1_More = 1'b1; $display(";A 2136");		//(= P1_P2_P1_More    0b1)) ;2136
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 2137");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b11101010)) ;2137
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2138");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2138
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2139");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2139
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2140");		//(= P1_P2_P1_Flush    0b0)) ;2140
                                    P1_P2_P1_More = 1'b0; $display(";A 2141");		//(= P1_P2_P1_More    0b0)) ;2141
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 2142");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b10110000)) ;2142
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2143");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2143
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2144");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2144
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2145");		//(= P1_P2_P1_Flush    0b0)) ;2145
                                    P1_P2_P1_More = 1'b0; $display(";A 2146");		//(= P1_P2_P1_More    0b0)) ;2146
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 2147");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b10111000)) ;2147
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 2148");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;2148
                                        P1_P2_P1_EAX <= #1 ((((P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 2150");		//(= P1_P2_P1_EAX    (bv-add (bv-add (bv-add (bv-mul P1_P2_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P2_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P2_P1_InstQueue 0  0b00000000000000000000000100000000)) P1_P2_P1_InstQueue 0 ))) ;2150
                                        P1_P2_P1_More = 1'b0; $display(";A 2151");		//(= P1_P2_P1_More    0b0)) ;2151
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2152");		//(= P1_P2_P1_Flush    0b0)) ;2152
                                        P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 2153");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;2153
                                        P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 2154");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;2154
                                    end
                                    else begin
                                        $display(";A 2149");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;2149
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2155");		//(= P1_P2_P1_Flush    0b0)) ;2155
                                        P1_P2_P1_More = 1'b1; $display(";A 2156");		//(= P1_P2_P1_More    0b1)) ;2156
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 2157");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b10111011)) ;2157
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 2158");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;2158
                                        P1_P2_P1_EBX <= #1 ((((P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P2_P1_InstQueue[((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 2160");		//(= P1_P2_P1_EBX    (bv-add (bv-add (bv-add (bv-mul P1_P2_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P2_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P2_P1_InstQueue 0  0b00000000000000000000000100000000)) P1_P2_P1_InstQueue 0 ))) ;2160
                                        P1_P2_P1_More = 1'b0; $display(";A 2161");		//(= P1_P2_P1_More    0b0)) ;2161
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2162");		//(= P1_P2_P1_Flush    0b0)) ;2162
                                        P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 2163");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;2163
                                        P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 2164");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;2164
                                    end
                                    else begin
                                        $display(";A 2159");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;2159
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2165");		//(= P1_P2_P1_Flush    0b0)) ;2165
                                        P1_P2_P1_More = 1'b1; $display(";A 2166");		//(= P1_P2_P1_More    0b1)) ;2166
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 2167");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b10001011)) ;2167
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2168");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2168
                                        if ((P1_P2_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 2170");		//(= (bool-to-bv (bv-slt P1_P2_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;2170
                                            P1_P2_P1_rEIP <= #1 (-P1_P2_P1_EBX); $display(";A 2172");		//(= P1_P2_P1_rEIP    (bv-neg P1_P2_P1_EBX ))) ;2172
                                        end
                                        else begin
                                            $display(";A 2171");		//(= (bool-to-bv (bv-slt P1_P2_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;2171
                                            P1_P2_P1_rEIP <= #1 P1_P2_P1_EBX; $display(";A 2173");		//(= P1_P2_P1_rEIP    P1_P2_P1_EBX )) ;2173
                                        end
                                        P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2174");		//(= P1_P2_P1_RequestPending    0b1)) ;2174
                                        P1_P2_P1_ReadRequest <= #1 1'b1; $display(";A 2175");		//(= P1_P2_P1_ReadRequest    0b1)) ;2175
                                        P1_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 2176");		//(= P1_P2_P1_MemoryFetch    0b1)) ;2176
                                        P1_P2_P1_CodeFetch <= #1 1'b0; $display(";A 2177");		//(= P1_P2_P1_CodeFetch    0b0)) ;2177
                                        if ((P1_P2_P1_READY_n == 1'b0)) begin
                                            $display(";A 2178");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2178
                                            P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2180");		//(= P1_P2_P1_RequestPending    0b0)) ;2180
                                            P1_P2_P1_uWord = (P1_P2_P1_Datai % 32'b00000000000000001000000000000000); $display(";A 2181");		//(= P1_P2_P1_uWord    (bv-smod P1_P2_P1_Datai  0b00000000000000001000000000000000))) ;2181
                                            if ((P1_P2_P1_StateBS16 == 1'b1)) begin
                                                $display(";A 2182");		//(= (bv-comp P1_P2_P1_StateBS16  0b1)   0b1)) ;2182
                                                P1_P2_P1_lWord = (P1_P2_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 2184");		//(= P1_P2_P1_lWord    (bv-smod P1_P2_P1_Datai  0b00000000000000010000000000000000))) ;2184
                                            end
                                            else begin
                                                $display(";A 2183");		//(= (bv-comp P1_P2_P1_StateBS16  0b1)   0b0)) ;2183
                                                P1_P2_P1_rEIP <= #1 (P1_P2_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 2185");		//(= P1_P2_P1_rEIP    (bv-add P1_P2_P1_rEIP  0b00000000000000000000000000000010))) ;2185
                                                P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2186");		//(= P1_P2_P1_RequestPending    0b1)) ;2186
                                                if ((P1_P2_P1_READY_n == 1'b0)) begin
                                                    $display(";A 2187");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2187
                                                    P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2189");		//(= P1_P2_P1_RequestPending    0b0)) ;2189
                                                    P1_P2_P1_lWord = (P1_P2_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 2190");		//(= P1_P2_P1_lWord    (bv-smod P1_P2_P1_Datai  0b00000000000000010000000000000000))) ;2190
                                                end
                                                else begin
                                                    $display(";A 2188");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2188
                                                end
                                            end
                                            if ((P1_P2_P1_READY_n == 1'b0)) begin
                                                $display(";A 2191");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2191
                                                P1_P2_P1_EAX <= #1 ((P1_P2_P1_uWord * 32'b00000000000000010000000000000000) + P1_P2_P1_lWord); $display(";A 2193");		//(= P1_P2_P1_EAX    (bv-add (bv-mul P1_P2_P1_uWord  0b00000000000000010000000000000000) P1_P2_P1_lWord ))) ;2193
                                                P1_P2_P1_More = 1'b0; $display(";A 2194");		//(= P1_P2_P1_More    0b0)) ;2194
                                                P1_P2_P1_Flush = 1'b0; $display(";A 2195");		//(= P1_P2_P1_Flush    0b0)) ;2195
                                                P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2196");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;2196
                                                P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2197");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2197
                                            end
                                            else begin
                                                $display(";A 2192");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2192
                                            end
                                        end
                                        else begin
                                            $display(";A 2179");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2179
                                        end
                                    end
                                    else begin
                                        $display(";A 2169");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2169
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2198");		//(= P1_P2_P1_Flush    0b0)) ;2198
                                        P1_P2_P1_More = 1'b1; $display(";A 2199");		//(= P1_P2_P1_More    0b1)) ;2199
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 2200");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b10001001)) ;2200
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2201");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2201
                                        if ((P1_P2_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 2203");		//(= (bool-to-bv (bv-slt P1_P2_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;2203
                                            P1_P2_P1_rEIP <= #1 P1_P2_P1_EBX; $display(";A 2205");		//(= P1_P2_P1_rEIP    P1_P2_P1_EBX )) ;2205
                                        end
                                        else begin
                                            $display(";A 2204");		//(= (bool-to-bv (bv-slt P1_P2_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;2204
                                            P1_P2_P1_rEIP <= #1 P1_P2_P1_EBX; $display(";A 2206");		//(= P1_P2_P1_rEIP    P1_P2_P1_EBX )) ;2206
                                        end
                                        P1_P2_P1_lWord = (P1_P2_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 2207");		//(= P1_P2_P1_lWord    (bv-smod P1_P2_P1_EAX  0b00000000000000010000000000000000))) ;2207
                                        P1_P2_P1_uWord = ((P1_P2_P1_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 2208");		//(= P1_P2_P1_uWord    (bv-smod (bv-sdiv P1_P2_P1_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;2208
                                        P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2209");		//(= P1_P2_P1_RequestPending    0b1)) ;2209
                                        P1_P2_P1_ReadRequest <= #1 1'b0; $display(";A 2210");		//(= P1_P2_P1_ReadRequest    0b0)) ;2210
                                        P1_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 2211");		//(= P1_P2_P1_MemoryFetch    0b1)) ;2211
                                        P1_P2_P1_CodeFetch <= #1 1'b0; $display(";A 2212");		//(= P1_P2_P1_CodeFetch    0b0)) ;2212
                                        if (((P1_P2_P1_State == 32'b00000000000000000000000000000010) | (P1_P2_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 2213");		//(= (bv-or (bv-comp P1_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P1_State  0b00000000000000000000000000000100))   0b1)) ;2213
                                            P1_P2_P1_Datao <= #1 ((P1_P2_P1_uWord * 32'b00000000000000010000000000000000) + P1_P2_P1_lWord); $display(";A 2215");		//(= P1_P2_P1_Datao    (bv-add (bv-mul P1_P2_P1_uWord  0b00000000000000010000000000000000) P1_P2_P1_lWord ))) ;2215
                                            if ((P1_P2_P1_READY_n == 1'b0)) begin
                                                $display(";A 2216");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2216
                                                P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2218");		//(= P1_P2_P1_RequestPending    0b0)) ;2218
                                                if ((P1_P2_P1_StateBS16 == 1'b0)) begin
                                                    $display(";A 2219");		//(= (bv-comp P1_P2_P1_StateBS16  0b0)   0b1)) ;2219
                                                    P1_P2_P1_rEIP <= #1 (P1_P2_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 2221");		//(= P1_P2_P1_rEIP    (bv-add P1_P2_P1_rEIP  0b00000000000000000000000000000010))) ;2221
                                                    P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2222");		//(= P1_P2_P1_RequestPending    0b1)) ;2222
                                                    P1_P2_P1_ReadRequest <= #1 1'b0; $display(";A 2223");		//(= P1_P2_P1_ReadRequest    0b0)) ;2223
                                                    P1_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 2224");		//(= P1_P2_P1_MemoryFetch    0b1)) ;2224
                                                    P1_P2_P1_CodeFetch <= #1 1'b0; $display(";A 2225");		//(= P1_P2_P1_CodeFetch    0b0)) ;2225
                                                    P1_P2_P1_State2 = 4'sb0110; $display(";A 2226");		//(= P1_P2_P1_State2    0b0110)) ;2226
                                                end
                                                else begin
                                                    $display(";A 2220");		//(= (bv-comp P1_P2_P1_StateBS16  0b0)   0b0)) ;2220
                                                end
                                                P1_P2_P1_More = 1'b0; $display(";A 2227");		//(= P1_P2_P1_More    0b0)) ;2227
                                                P1_P2_P1_Flush = 1'b0; $display(";A 2228");		//(= P1_P2_P1_Flush    0b0)) ;2228
                                                P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2229");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;2229
                                                P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2230");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2230
                                            end
                                            else begin
                                                $display(";A 2217");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2217
                                            end
                                        end
                                        else begin
                                            $display(";A 2214");		//(= (bv-or (bv-comp P1_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P1_State  0b00000000000000000000000000000100))   0b0)) ;2214
                                        end
                                    end
                                    else begin
                                        $display(";A 2202");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2202
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2231");		//(= P1_P2_P1_Flush    0b0)) ;2231
                                        P1_P2_P1_More = 1'b1; $display(";A 2232");		//(= P1_P2_P1_More    0b1)) ;2232
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 2233");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b11100100)) ;2233
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2234");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2234
                                        P1_P2_P1_rEIP <= #1 (P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 2236");		//(= P1_P2_P1_rEIP    (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;2236
                                        P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2237");		//(= P1_P2_P1_RequestPending    0b1)) ;2237
                                        P1_P2_P1_ReadRequest <= #1 1'b1; $display(";A 2238");		//(= P1_P2_P1_ReadRequest    0b1)) ;2238
                                        P1_P2_P1_MemoryFetch <= #1 1'b0; $display(";A 2239");		//(= P1_P2_P1_MemoryFetch    0b0)) ;2239
                                        P1_P2_P1_CodeFetch <= #1 1'b0; $display(";A 2240");		//(= P1_P2_P1_CodeFetch    0b0)) ;2240
                                        if ((P1_P2_P1_READY_n == 1'b0)) begin
                                            $display(";A 2241");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2241
                                            P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2243");		//(= P1_P2_P1_RequestPending    0b0)) ;2243
                                            P1_P2_P1_EAX <= #1 P1_P2_P1_Datai; $display(";A 2244");		//(= P1_P2_P1_EAX    P1_P2_P1_Datai )) ;2244
                                            P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2245");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;2245
                                            P1_P2_P1_InstQueueRd_Addr = (P1_P2_P1_InstQueueRd_Addr + 5'b00010); $display(";A 2246");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-add P1_P2_P1_InstQueueRd_Addr  0b00010))) ;2246
                                            P1_P2_P1_Flush = 1'b0; $display(";A 2247");		//(= P1_P2_P1_Flush    0b0)) ;2247
                                            P1_P2_P1_More = 1'b0; $display(";A 2248");		//(= P1_P2_P1_More    0b0)) ;2248
                                        end
                                        else begin
                                            $display(";A 2242");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2242
                                        end
                                    end
                                    else begin
                                        $display(";A 2235");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2235
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2249");		//(= P1_P2_P1_Flush    0b0)) ;2249
                                        P1_P2_P1_More = 1'b1; $display(";A 2250");		//(= P1_P2_P1_More    0b1)) ;2250
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 2251");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b11100110)) ;2251
                                    if (((P1_P2_P1_InstQueueWr_Addr - P1_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2252");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2252
                                        P1_P2_P1_rEIP <= #1 (P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 2254");		//(= P1_P2_P1_rEIP    (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;2254
                                        P1_P2_P1_RequestPending <= #1 1'b1; $display(";A 2255");		//(= P1_P2_P1_RequestPending    0b1)) ;2255
                                        P1_P2_P1_ReadRequest <= #1 1'b0; $display(";A 2256");		//(= P1_P2_P1_ReadRequest    0b0)) ;2256
                                        P1_P2_P1_MemoryFetch <= #1 1'b0; $display(";A 2257");		//(= P1_P2_P1_MemoryFetch    0b0)) ;2257
                                        P1_P2_P1_CodeFetch <= #1 1'b0; $display(";A 2258");		//(= P1_P2_P1_CodeFetch    0b0)) ;2258
                                        if (((P1_P2_P1_State == 32'b00000000000000000000000000000010) | (P1_P2_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 2259");		//(= (bv-or (bv-comp P1_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P1_State  0b00000000000000000000000000000100))   0b1)) ;2259
                                            P1_P2_P1_fWord = (P1_P2_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 2261");		//(= P1_P2_P1_fWord    (bv-smod P1_P2_P1_EAX  0b00000000000000010000000000000000))) ;2261
                                            P1_P2_P1_Datao <= #1 P1_P2_P1_fWord; $display(";A 2262");		//(= P1_P2_P1_Datao    P1_P2_P1_fWord )) ;2262
                                            if ((P1_P2_P1_READY_n == 1'b0)) begin
                                                $display(";A 2263");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2263
                                                P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2265");		//(= P1_P2_P1_RequestPending    0b0)) ;2265
                                                P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2266");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;2266
                                                P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2267");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2267
                                                P1_P2_P1_Flush = 1'b0; $display(";A 2268");		//(= P1_P2_P1_Flush    0b0)) ;2268
                                                P1_P2_P1_More = 1'b0; $display(";A 2269");		//(= P1_P2_P1_More    0b0)) ;2269
                                            end
                                            else begin
                                                $display(";A 2264");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2264
                                            end
                                        end
                                        else begin
                                            $display(";A 2260");		//(= (bv-or (bv-comp P1_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P1_State  0b00000000000000000000000000000100))   0b0)) ;2260
                                        end
                                    end
                                    else begin
                                        $display(";A 2253");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P1_InstQueueWr_Addr  P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2253
                                        P1_P2_P1_Flush = 1'b0; $display(";A 2270");		//(= P1_P2_P1_Flush    0b0)) ;2270
                                        P1_P2_P1_More = 1'b1; $display(";A 2271");		//(= P1_P2_P1_More    0b1)) ;2271
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 2272");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b00000100)) ;2272
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2273");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2273
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2274");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2274
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2275");		//(= P1_P2_P1_Flush    0b0)) ;2275
                                    P1_P2_P1_More = 1'b0; $display(";A 2276");		//(= P1_P2_P1_More    0b0)) ;2276
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 2277");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b00000101)) ;2277
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2278");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2278
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2279");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2279
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2280");		//(= P1_P2_P1_Flush    0b0)) ;2280
                                    P1_P2_P1_More = 1'b0; $display(";A 2281");		//(= P1_P2_P1_More    0b0)) ;2281
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 2282");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b11010000)) ;2282
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2283");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;2283
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2284");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2284
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2285");		//(= P1_P2_P1_Flush    0b0)) ;2285
                                    P1_P2_P1_More = 1'b0; $display(";A 2286");		//(= P1_P2_P1_More    0b0)) ;2286
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 2287");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b11000000)) ;2287
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2288");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;2288
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2289");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2289
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2290");		//(= P1_P2_P1_Flush    0b0)) ;2290
                                    P1_P2_P1_More = 1'b0; $display(";A 2291");		//(= P1_P2_P1_More    0b0)) ;2291
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 2292");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b01000000)) ;2292
                                    P1_P2_P1_EAX <= #1 (P1_P2_P1_EAX + 32'sb00000000000000000000000000000001); $display(";A 2293");		//(= P1_P2_P1_EAX    (bv-add P1_P2_P1_EAX  0b00000000000000000000000000000001))) ;2293
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2294");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2294
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2295");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2295
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2296");		//(= P1_P2_P1_Flush    0b0)) ;2296
                                    P1_P2_P1_More = 1'b0; $display(";A 2297");		//(= P1_P2_P1_More    0b0)) ;2297
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 2298");		//(= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr )   0b01000011)) ;2298
                                    P1_P2_P1_EBX <= #1 (P1_P2_P1_EBX + 32'sb00000000000000000000000000000001); $display(";A 2299");		//(= P1_P2_P1_EBX    (bv-add P1_P2_P1_EBX  0b00000000000000000000000000000001))) ;2299
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2300");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2300
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2301");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2301
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2302");		//(= P1_P2_P1_Flush    0b0)) ;2302
                                    P1_P2_P1_More = 1'b0; $display(";A 2303");		//(= P1_P2_P1_More    0b0)) ;2303
                                end
                            default:
                                begin
                                    $display(";A 2304");		//(= (and (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b10010000) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b01100110) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b11101011) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b11101001) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b11101010) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b10110000) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b10111000) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b10111011) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b10001011) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b10001001) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b11100100) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b11100110) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b00000100) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b00000101) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b11010000) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b11000000) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b01000000) (/= ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ) 0b01000011))   true)) ;2304
                                    P1_P2_P1_InstAddrPointer = (P1_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2305");		//(= P1_P2_P1_InstAddrPointer    (bv-add P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;2305
                                    P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2306");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2306
                                    P1_P2_P1_Flush = 1'b0; $display(";A 2307");		//(= P1_P2_P1_Flush    0b0)) ;2307
                                    P1_P2_P1_More = 1'b0; $display(";A 2308");		//(= P1_P2_P1_More    0b0)) ;2308
                                end
                        endcase
                        if (((~(P1_P2_P1_InstQueueRd_Addr < P1_P2_P1_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P1_P2_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P1_P2_P1_Flush) | P1_P2_P1_More))) begin
                            $display(";A 2309");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P2_P1_InstQueueRd_Addr  P1_P2_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P2_P1_Flush ) P1_P2_P1_More ))   0b1)) ;2309
                            P1_P2_P1_State2 = 4'sb0111; $display(";A 2311");		//(= P1_P2_P1_State2    0b0111)) ;2311
                        end
                        else begin
                            $display(";A 2310");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P2_P1_InstQueueRd_Addr  P1_P2_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P2_P1_Flush ) P1_P2_P1_More ))   0b0)) ;2310
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 2312");		//(= P1_P2_P1_State2    0b0110)) ;2312
                        P1_P2_P1_Datao <= #1 ((P1_P2_P1_uWord * 32'b00000000000000010000000000000000) + P1_P2_P1_lWord); $display(";A 2313");		//(= P1_P2_P1_Datao    (bv-add (bv-mul P1_P2_P1_uWord  0b00000000000000010000000000000000) P1_P2_P1_lWord ))) ;2313
                        if ((P1_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 2314");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b1)) ;2314
                            P1_P2_P1_RequestPending <= #1 1'b0; $display(";A 2316");		//(= P1_P2_P1_RequestPending    0b0)) ;2316
                            P1_P2_P1_State2 = 4'sb0101; $display(";A 2317");		//(= P1_P2_P1_State2    0b0101)) ;2317
                        end
                        else begin
                            $display(";A 2315");		//(= (bv-comp P1_P2_P1_READY_n  0b0)   0b0)) ;2315
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 2318");		//(= P1_P2_P1_State2    0b0111)) ;2318
                        if (P1_P2_P1_Flush) begin
                            $display(";A 2319");		//(= P1_P2_P1_Flush    0b1)) ;2319
                            P1_P2_P1_InstQueueRd_Addr = 5'sb00001; $display(";A 2321");		//(= P1_P2_P1_InstQueueRd_Addr    0b00001)) ;2321
                            P1_P2_P1_InstQueueWr_Addr = 5'sb00001; $display(";A 2322");		//(= P1_P2_P1_InstQueueWr_Addr    0b00001)) ;2322
                            if ((P1_P2_P1_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 2323");		//(= (bool-to-bv (bv-slt P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;2323
                                P1_P2_P1_fWord = (-P1_P2_P1_InstAddrPointer); $display(";A 2325");		//(= P1_P2_P1_fWord    (bv-neg P1_P2_P1_InstAddrPointer ))) ;2325
                            end
                            else begin
                                $display(";A 2324");		//(= (bool-to-bv (bv-slt P1_P2_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;2324
                                P1_P2_P1_fWord = P1_P2_P1_InstAddrPointer; $display(";A 2326");		//(= P1_P2_P1_fWord    P1_P2_P1_InstAddrPointer )) ;2326
                            end
                            if (((P1_P2_P1_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 2327");		//(= (bv-comp (bv-smod P1_P2_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;2327
                                P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + (P1_P2_P1_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 2329");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  (bv-smod P1_P2_P1_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;2329
                            end
                            else begin
                                $display(";A 2328");		//(= (bv-comp (bv-smod P1_P2_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;2328
                            end
                        end
                        else begin
                            $display(";A 2320");		//(= P1_P2_P1_Flush    0b0)) ;2320
                        end
                        if (((32'b00000000000000000000000000001111 - P1_P2_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 2330");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;2330
                            P1_P2_P1_State2 = 4'sb1000; $display(";A 2332");		//(= P1_P2_P1_State2    0b1000)) ;2332
                            P1_P2_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 2333");		//(= P1_P2_P1_InstQueueWr_Addr    0b00000)) ;2333
                        end
                        else begin
                            $display(";A 2331");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;2331
                            P1_P2_P1_State2 = 4'sb1001; $display(";A 2334");		//(= P1_P2_P1_State2    0b1001)) ;2334
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 2335");		//(= P1_P2_P1_State2    0b1000)) ;2335
                        if ((P1_P2_P1_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 2336");		//(= (bool-to-bv (bv-le P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;2336
                            P1_P2_P1_InstQueue[P1_P2_P1_InstQueueWr_Addr] = P1_P2_P1_InstQueue[P1_P2_P1_InstQueueRd_Addr]; $display(";A 2338");		//(= P1_P2_P1_InstQueue    ( P1_P2_P1_InstQueue P1_P2_P1_InstQueueRd_Addr ))) ;2338
                            P1_P2_P1_InstQueueRd_Addr = ((P1_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2339");		//(= P1_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2339
                            P1_P2_P1_InstQueueWr_Addr = ((P1_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2340");		//(= P1_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2340
                            P1_P2_P1_State2 = 4'sb1000; $display(";A 2341");		//(= P1_P2_P1_State2    0b1000)) ;2341
                        end
                        else begin
                            $display(";A 2337");		//(= (bool-to-bv (bv-le P1_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;2337
                            P1_P2_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 2342");		//(= P1_P2_P1_InstQueueRd_Addr    0b00000)) ;2342
                            P1_P2_P1_State2 = 4'sb1001; $display(";A 2343");		//(= P1_P2_P1_State2    0b1001)) ;2343
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 2344");		//(= P1_P2_P1_State2    0b1001)) ;2344
                        P1_P2_P1_rEIP <= #1 P1_P2_P1_PhyAddrPointer; $display(";A 2345");		//(= P1_P2_P1_rEIP    P1_P2_P1_PhyAddrPointer )) ;2345
                        P1_P2_P1_State2 = 4'sb0001; $display(";A 2346");		//(= P1_P2_P1_State2    0b0001)) ;2346
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:3398
    always @(posedge P1_P2_P1_RESET or posedge P1_P2_P1_CLOCK) begin
        if ((P1_P2_P1_RESET == 1'b1)) begin
            $display(";A 2347");		//(= (bv-comp P1_P2_P1_RESET  0b1)   0b1)) ;2347
            P1_P2_P1_ByteEnable <= #1 4'b0000; $display(";A 2349");		//(= P1_P2_P1_ByteEnable    0b0000)) ;2349
            P1_P2_P1_NonAligned <= #1 1'b0; $display(";A 2350");		//(= P1_P2_P1_NonAligned    0b0)) ;2350
        end
        else begin
            $display(";A 2348");		//(= (bv-comp P1_P2_P1_RESET  0b1)   0b0)) ;2348
            case (P1_P2_P1_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 2351");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000000)) ;2351
                        case ((P1_P2_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 2352");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;2352
                                    P1_P2_P1_ByteEnable <= #1 4'b1110; $display(";A 2353");		//(= P1_P2_P1_ByteEnable    0b1110)) ;2353
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 2354");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;2354
                                    P1_P2_P1_ByteEnable <= #1 4'b1101; $display(";A 2355");		//(= P1_P2_P1_ByteEnable    0b1101)) ;2355
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 2356");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;2356
                                    P1_P2_P1_ByteEnable <= #1 4'b1011; $display(";A 2357");		//(= P1_P2_P1_ByteEnable    0b1011)) ;2357
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 2358");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;2358
                                    P1_P2_P1_ByteEnable <= #1 4'b0111; $display(";A 2359");		//(= P1_P2_P1_ByteEnable    0b0111)) ;2359
                                end
                            default:
                                begin
                                    $display(";A 2360");		//(= (and (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;2360
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 2361");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000001)) ;2361
                        case ((P1_P2_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 2362");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;2362
                                    P1_P2_P1_ByteEnable <= #1 4'b1100; $display(";A 2363");		//(= P1_P2_P1_ByteEnable    0b1100)) ;2363
                                    P1_P2_P1_NonAligned <= #1 1'b0; $display(";A 2364");		//(= P1_P2_P1_NonAligned    0b0)) ;2364
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 2365");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;2365
                                    P1_P2_P1_ByteEnable <= #1 4'b1001; $display(";A 2366");		//(= P1_P2_P1_ByteEnable    0b1001)) ;2366
                                    P1_P2_P1_NonAligned <= #1 1'b0; $display(";A 2367");		//(= P1_P2_P1_NonAligned    0b0)) ;2367
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 2368");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;2368
                                    P1_P2_P1_ByteEnable <= #1 4'b0011; $display(";A 2369");		//(= P1_P2_P1_ByteEnable    0b0011)) ;2369
                                    P1_P2_P1_NonAligned <= #1 1'b0; $display(";A 2370");		//(= P1_P2_P1_NonAligned    0b0)) ;2370
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 2371");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;2371
                                    P1_P2_P1_ByteEnable <= #1 4'b0111; $display(";A 2372");		//(= P1_P2_P1_ByteEnable    0b0111)) ;2372
                                    P1_P2_P1_NonAligned <= #1 1'b1; $display(";A 2373");		//(= P1_P2_P1_NonAligned    0b1)) ;2373
                                end
                            default:
                                begin
                                    $display(";A 2374");		//(= (and (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;2374
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 2375");		//(= P1_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;2375
                        case ((P1_P2_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 2376");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;2376
                                    P1_P2_P1_ByteEnable <= #1 4'b0000; $display(";A 2377");		//(= P1_P2_P1_ByteEnable    0b0000)) ;2377
                                    P1_P2_P1_NonAligned <= #1 1'b0; $display(";A 2378");		//(= P1_P2_P1_NonAligned    0b0)) ;2378
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 2379");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;2379
                                    P1_P2_P1_ByteEnable <= #1 4'b0001; $display(";A 2380");		//(= P1_P2_P1_ByteEnable    0b0001)) ;2380
                                    P1_P2_P1_NonAligned <= #1 1'b1; $display(";A 2381");		//(= P1_P2_P1_NonAligned    0b1)) ;2381
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 2382");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;2382
                                    P1_P2_P1_NonAligned <= #1 1'b1; $display(";A 2383");		//(= P1_P2_P1_NonAligned    0b1)) ;2383
                                    P1_P2_P1_ByteEnable <= #1 4'b0011; $display(";A 2384");		//(= P1_P2_P1_ByteEnable    0b0011)) ;2384
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 2385");		//(= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;2385
                                    P1_P2_P1_NonAligned <= #1 1'b1; $display(";A 2386");		//(= P1_P2_P1_NonAligned    0b1)) ;2386
                                    P1_P2_P1_ByteEnable <= #1 4'b0111; $display(";A 2387");		//(= P1_P2_P1_ByteEnable    0b0111)) ;2387
                                end
                            default:
                                begin
                                    $display(";A 2388");		//(= (and (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;2388
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 2389");		//(= (and (/= P1_P2_P1_DataWidth  0b00000000000000000000000000000000) (/= P1_P2_P1_DataWidth  0b00000000000000000000000000000001) (/= P1_P2_P1_DataWidth  0b00000000000000000000000000000010))   true)) ;2389
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:3586
    always @(posedge P1_P2_P2_RESET or posedge P1_P2_P2_CLOCK) begin
        if ((P1_P2_P2_RESET == 1'b1)) begin
            $display(";A 2390");		//(= (bv-comp P1_P2_P2_RESET  0b1)   0b1)) ;2390
            P1_P2_P2_BE_n <= #1 4'b0000; $display(";A 2392");		//(= P1_P2_P2_BE_n    0b0000)) ;2392
            P1_P2_P2_Address <= #1 30'sb000000000000000000000000000000; $display(";A 2393");		//(= P1_P2_P2_Address    0b000000000000000000000000000000)) ;2393
            P1_P2_P2_W_R_n <= #1 1'b0; $display(";A 2394");		//(= P1_P2_P2_W_R_n    0b0)) ;2394
            P1_P2_P2_D_C_n <= #1 1'b0; $display(";A 2395");		//(= P1_P2_P2_D_C_n    0b0)) ;2395
            P1_P2_P2_M_IO_n <= #1 1'b0; $display(";A 2396");		//(= P1_P2_P2_M_IO_n    0b0)) ;2396
            P1_P2_P2_ADS_n <= #1 1'b0; $display(";A 2397");		//(= P1_P2_P2_ADS_n    0b0)) ;2397
            P1_P2_P2_State <= #1 3'sb000; $display(";A 2398");		//(= P1_P2_P2_State    0b000)) ;2398
            P1_P2_P2_StateNA <= #1 1'b0; $display(";A 2399");		//(= P1_P2_P2_StateNA    0b0)) ;2399
            P1_P2_P2_StateBS16 <= #1 1'b0; $display(";A 2400");		//(= P1_P2_P2_StateBS16    0b0)) ;2400
            P1_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 2401");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000000)) ;2401
        end
        else begin
            $display(";A 2391");		//(= (bv-comp P1_P2_P2_RESET  0b1)   0b0)) ;2391
            case (P1_P2_P2_State)
                3'b000 :
                    begin
                        $display(";A 2402");		//(= P1_P2_P2_State    0b000)) ;2402
                        P1_P2_P2_D_C_n <= #1 1'b1; $display(";A 2403");		//(= P1_P2_P2_D_C_n    0b1)) ;2403
                        P1_P2_P2_ADS_n <= #1 1'b1; $display(";A 2404");		//(= P1_P2_P2_ADS_n    0b1)) ;2404
                        P1_P2_P2_State <= #1 3'sb001; $display(";A 2405");		//(= P1_P2_P2_State    0b001)) ;2405
                        P1_P2_P2_StateNA <= #1 1'b1; $display(";A 2406");		//(= P1_P2_P2_StateNA    0b1)) ;2406
                        P1_P2_P2_StateBS16 <= #1 1'b1; $display(";A 2407");		//(= P1_P2_P2_StateBS16    0b1)) ;2407
                        P1_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 2408");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;2408
                        P1_P2_P2_State <= #1 3'sb001; $display(";A 2409");		//(= P1_P2_P2_State    0b001)) ;2409
                    end
                3'b001 :
                    begin
                        $display(";A 2410");		//(= P1_P2_P2_State    0b001)) ;2410
                        if ((P1_P2_P2_RequestPending == 1'b1)) begin
                            $display(";A 2411");		//(= (bv-comp P1_P2_P2_RequestPending  0b1)   0b1)) ;2411
                            P1_P2_P2_State <= #1 3'sb010; $display(";A 2413");		//(= P1_P2_P2_State    0b010)) ;2413
                        end
                        else begin
                            $display(";A 2412");		//(= (bv-comp P1_P2_P2_RequestPending  0b1)   0b0)) ;2412
                            if ((P1_P2_P2_HOLD == 1'b1)) begin
                                $display(";A 2414");		//(= (bv-comp P1_P2_P2_HOLD  0b1)   0b1)) ;2414
                                P1_P2_P2_State <= #1 3'sb101; $display(";A 2416");		//(= P1_P2_P2_State    0b101)) ;2416
                            end
                            else begin
                                $display(";A 2415");		//(= (bv-comp P1_P2_P2_HOLD  0b1)   0b0)) ;2415
                                P1_P2_P2_State <= #1 3'sb001; $display(";A 2417");		//(= P1_P2_P2_State    0b001)) ;2417
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 2418");		//(= P1_P2_P2_State    0b010)) ;2418
                        P1_P2_P2_Address <= #1 ((P1_P2_P2_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 2419");		//(= P1_P2_P2_Address    (bv-smod (bv-sdiv P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;2419
                        P1_P2_P2_BE_n <= #1 P1_P2_P2_ByteEnable; $display(";A 2420");		//(= P1_P2_P2_BE_n    P1_P2_P2_ByteEnable )) ;2420
                        P1_P2_P2_M_IO_n <= #1 P1_P2_P2_MemoryFetch; $display(";A 2421");		//(= P1_P2_P2_M_IO_n    P1_P2_P2_MemoryFetch )) ;2421
                        if ((P1_P2_P2_ReadRequest == 1'b1)) begin
                            $display(";A 2422");		//(= (bv-comp P1_P2_P2_ReadRequest  0b1)   0b1)) ;2422
                            P1_P2_P2_W_R_n <= #1 1'b0; $display(";A 2424");		//(= P1_P2_P2_W_R_n    0b0)) ;2424
                        end
                        else begin
                            $display(";A 2423");		//(= (bv-comp P1_P2_P2_ReadRequest  0b1)   0b0)) ;2423
                            P1_P2_P2_W_R_n <= #1 1'b1; $display(";A 2425");		//(= P1_P2_P2_W_R_n    0b1)) ;2425
                        end
                        if ((P1_P2_P2_CodeFetch == 1'b1)) begin
                            $display(";A 2426");		//(= (bv-comp P1_P2_P2_CodeFetch  0b1)   0b1)) ;2426
                            P1_P2_P2_D_C_n <= #1 1'b0; $display(";A 2428");		//(= P1_P2_P2_D_C_n    0b0)) ;2428
                        end
                        else begin
                            $display(";A 2427");		//(= (bv-comp P1_P2_P2_CodeFetch  0b1)   0b0)) ;2427
                            P1_P2_P2_D_C_n <= #1 1'b1; $display(";A 2429");		//(= P1_P2_P2_D_C_n    0b1)) ;2429
                        end
                        P1_P2_P2_ADS_n <= #1 1'b0; $display(";A 2430");		//(= P1_P2_P2_ADS_n    0b0)) ;2430
                        P1_P2_P2_State <= #1 3'sb011; $display(";A 2431");		//(= P1_P2_P2_State    0b011)) ;2431
                    end
                3'b011 :
                    begin
                        $display(";A 2432");		//(= P1_P2_P2_State    0b011)) ;2432
                        if ((((P1_P2_P2_READY_n == 1'b0) & (P1_P2_P2_HOLD == 1'b0)) & (P1_P2_P2_RequestPending == 1'b1))) begin
                            $display(";A 2433");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b1))   0b1)) ;2433
                            P1_P2_P2_State <= #1 3'sb010; $display(";A 2435");		//(= P1_P2_P2_State    0b010)) ;2435
                        end
                        else begin
                            $display(";A 2434");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b1))   0b0)) ;2434
                            if (((P1_P2_P2_READY_n == 1'b1) & (P1_P2_P2_NA_n == 1'b1))) begin
                                $display(";A 2436");		//(= (bv-and (bv-comp P1_P2_P2_READY_n  0b1) (bv-comp P1_P2_P2_NA_n  0b1))   0b1)) ;2436
                            end
                            else begin
                                $display(";A 2437");		//(= (bv-and (bv-comp P1_P2_P2_READY_n  0b1) (bv-comp P1_P2_P2_NA_n  0b1))   0b0)) ;2437
                                if ((((P1_P2_P2_RequestPending == 1'b1) | (P1_P2_P2_HOLD == 1'b1)) & ((P1_P2_P2_READY_n == 1'b1) & (P1_P2_P2_NA_n == 1'b0)))) begin
                                    $display(";A 2438");		//(= (bv-and (bv-or (bv-comp P1_P2_P2_RequestPending  0b1) (bv-comp P1_P2_P2_HOLD  0b1)) (bv-and (bv-comp P1_P2_P2_READY_n  0b1) (bv-comp P1_P2_P2_NA_n  0b0)))   0b1)) ;2438
                                    P1_P2_P2_State <= #1 3'sb111; $display(";A 2440");		//(= P1_P2_P2_State    0b111)) ;2440
                                end
                                else begin
                                    $display(";A 2439");		//(= (bv-and (bv-or (bv-comp P1_P2_P2_RequestPending  0b1) (bv-comp P1_P2_P2_HOLD  0b1)) (bv-and (bv-comp P1_P2_P2_READY_n  0b1) (bv-comp P1_P2_P2_NA_n  0b0)))   0b0)) ;2439
                                    if (((((P1_P2_P2_RequestPending == 1'b1) & (P1_P2_P2_HOLD == 1'b0)) & (P1_P2_P2_READY_n == 1'b1)) & (P1_P2_P2_NA_n == 1'b0))) begin
                                        $display(";A 2441");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P2_P2_RequestPending  0b1) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_READY_n  0b1)) (bv-comp P1_P2_P2_NA_n  0b0))   0b1)) ;2441
                                        P1_P2_P2_State <= #1 3'sb110; $display(";A 2443");		//(= P1_P2_P2_State    0b110)) ;2443
                                    end
                                    else begin
                                        $display(";A 2442");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P2_P2_RequestPending  0b1) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_READY_n  0b1)) (bv-comp P1_P2_P2_NA_n  0b0))   0b0)) ;2442
                                        if ((((P1_P2_P2_RequestPending == 1'b0) & (P1_P2_P2_HOLD == 1'b0)) & (P1_P2_P2_READY_n == 1'b0))) begin
                                            $display(";A 2444");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_RequestPending  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_READY_n  0b0))   0b1)) ;2444
                                            P1_P2_P2_State <= #1 3'sb001; $display(";A 2446");		//(= P1_P2_P2_State    0b001)) ;2446
                                        end
                                        else begin
                                            $display(";A 2445");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_RequestPending  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_READY_n  0b0))   0b0)) ;2445
                                            if (((P1_P2_P2_HOLD == 1'b1) & (P1_P2_P2_READY_n == 1'b1))) begin
                                                $display(";A 2447");		//(= (bv-and (bv-comp P1_P2_P2_HOLD  0b1) (bv-comp P1_P2_P2_READY_n  0b1))   0b1)) ;2447
                                                P1_P2_P2_State <= #1 3'sb101; $display(";A 2449");		//(= P1_P2_P2_State    0b101)) ;2449
                                            end
                                            else begin
                                                $display(";A 2448");		//(= (bv-and (bv-comp P1_P2_P2_HOLD  0b1) (bv-comp P1_P2_P2_READY_n  0b1))   0b0)) ;2448
                                                P1_P2_P2_State <= #1 3'sb011; $display(";A 2450");		//(= P1_P2_P2_State    0b011)) ;2450
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P1_P2_P2_StateBS16 <= #1 P1_P2_P2_BS16_n; $display(";A 2451");		//(= P1_P2_P2_StateBS16    P1_P2_P2_BS16_n )) ;2451
                        if ((P1_P2_P2_BS16_n == 1'b0)) begin
                            $display(";A 2452");		//(= (bv-comp P1_P2_P2_BS16_n  0b0)   0b1)) ;2452
                            P1_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 2454");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000001)) ;2454
                        end
                        else begin
                            $display(";A 2453");		//(= (bv-comp P1_P2_P2_BS16_n  0b0)   0b0)) ;2453
                            P1_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 2455");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;2455
                        end
                        P1_P2_P2_StateNA <= #1 P1_P2_P2_NA_n; $display(";A 2456");		//(= P1_P2_P2_StateNA    P1_P2_P2_NA_n )) ;2456
                        P1_P2_P2_ADS_n <= #1 1'b1; $display(";A 2457");		//(= P1_P2_P2_ADS_n    0b1)) ;2457
                    end
                3'b100 :
                    begin
                        $display(";A 2458");		//(= P1_P2_P2_State    0b100)) ;2458
                        if ((((P1_P2_P2_NA_n == 1'b0) & (P1_P2_P2_HOLD == 1'b0)) & (P1_P2_P2_RequestPending == 1'b1))) begin
                            $display(";A 2459");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_NA_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b1))   0b1)) ;2459
                            P1_P2_P2_State <= #1 3'sb110; $display(";A 2461");		//(= P1_P2_P2_State    0b110)) ;2461
                        end
                        else begin
                            $display(";A 2460");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_NA_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b1))   0b0)) ;2460
                            if (((P1_P2_P2_NA_n == 1'b0) & ((P1_P2_P2_HOLD == 1'b1) | (P1_P2_P2_RequestPending == 1'b0)))) begin
                                $display(";A 2462");		//(= (bv-and (bv-comp P1_P2_P2_NA_n  0b0) (bv-or (bv-comp P1_P2_P2_HOLD  0b1) (bv-comp P1_P2_P2_RequestPending  0b0)))   0b1)) ;2462
                                P1_P2_P2_State <= #1 3'sb111; $display(";A 2464");		//(= P1_P2_P2_State    0b111)) ;2464
                            end
                            else begin
                                $display(";A 2463");		//(= (bv-and (bv-comp P1_P2_P2_NA_n  0b0) (bv-or (bv-comp P1_P2_P2_HOLD  0b1) (bv-comp P1_P2_P2_RequestPending  0b0)))   0b0)) ;2463
                                if ((P1_P2_P2_NA_n == 1'b1)) begin
                                    $display(";A 2465");		//(= (bv-comp P1_P2_P2_NA_n  0b1)   0b1)) ;2465
                                    P1_P2_P2_State <= #1 3'sb011; $display(";A 2467");		//(= P1_P2_P2_State    0b011)) ;2467
                                end
                                else begin
                                    $display(";A 2466");		//(= (bv-comp P1_P2_P2_NA_n  0b1)   0b0)) ;2466
                                    P1_P2_P2_State <= #1 3'sb100; $display(";A 2468");		//(= P1_P2_P2_State    0b100)) ;2468
                                end
                            end
                        end
                        P1_P2_P2_StateBS16 <= #1 P1_P2_P2_BS16_n; $display(";A 2469");		//(= P1_P2_P2_StateBS16    P1_P2_P2_BS16_n )) ;2469
                        if ((P1_P2_P2_BS16_n == 1'b0)) begin
                            $display(";A 2470");		//(= (bv-comp P1_P2_P2_BS16_n  0b0)   0b1)) ;2470
                            P1_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 2472");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000001)) ;2472
                        end
                        else begin
                            $display(";A 2471");		//(= (bv-comp P1_P2_P2_BS16_n  0b0)   0b0)) ;2471
                            P1_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 2473");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;2473
                        end
                        P1_P2_P2_StateNA <= #1 P1_P2_P2_NA_n; $display(";A 2474");		//(= P1_P2_P2_StateNA    P1_P2_P2_NA_n )) ;2474
                        P1_P2_P2_ADS_n <= #1 1'b1; $display(";A 2475");		//(= P1_P2_P2_ADS_n    0b1)) ;2475
                    end
                3'b101 :
                    begin
                        $display(";A 2476");		//(= P1_P2_P2_State    0b101)) ;2476
                        if (((P1_P2_P2_HOLD == 1'b0) & (P1_P2_P2_RequestPending == 1'b1))) begin
                            $display(";A 2477");		//(= (bv-and (bv-comp P1_P2_P2_HOLD  0b0) (bv-comp P1_P2_P2_RequestPending  0b1))   0b1)) ;2477
                            P1_P2_P2_State <= #1 3'sb010; $display(";A 2479");		//(= P1_P2_P2_State    0b010)) ;2479
                        end
                        else begin
                            $display(";A 2478");		//(= (bv-and (bv-comp P1_P2_P2_HOLD  0b0) (bv-comp P1_P2_P2_RequestPending  0b1))   0b0)) ;2478
                            if (((P1_P2_P2_HOLD == 1'b0) & (P1_P2_P2_RequestPending == 1'b0))) begin
                                $display(";A 2480");		//(= (bv-and (bv-comp P1_P2_P2_HOLD  0b0) (bv-comp P1_P2_P2_RequestPending  0b0))   0b1)) ;2480
                                P1_P2_P2_State <= #1 3'sb001; $display(";A 2482");		//(= P1_P2_P2_State    0b001)) ;2482
                            end
                            else begin
                                $display(";A 2481");		//(= (bv-and (bv-comp P1_P2_P2_HOLD  0b0) (bv-comp P1_P2_P2_RequestPending  0b0))   0b0)) ;2481
                                P1_P2_P2_State <= #1 3'sb101; $display(";A 2483");		//(= P1_P2_P2_State    0b101)) ;2483
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 2484");		//(= P1_P2_P2_State    0b110)) ;2484
                        P1_P2_P2_Address <= #1 ((P1_P2_P2_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 2485");		//(= P1_P2_P2_Address    (bv-smod (bv-sdiv P1_P2_P2_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;2485
                        P1_P2_P2_BE_n <= #1 P1_P2_P2_ByteEnable; $display(";A 2486");		//(= P1_P2_P2_BE_n    P1_P2_P2_ByteEnable )) ;2486
                        P1_P2_P2_M_IO_n <= #1 P1_P2_P2_MemoryFetch; $display(";A 2487");		//(= P1_P2_P2_M_IO_n    P1_P2_P2_MemoryFetch )) ;2487
                        if ((P1_P2_P2_ReadRequest == 1'b1)) begin
                            $display(";A 2488");		//(= (bv-comp P1_P2_P2_ReadRequest  0b1)   0b1)) ;2488
                            P1_P2_P2_W_R_n <= #1 1'b0; $display(";A 2490");		//(= P1_P2_P2_W_R_n    0b0)) ;2490
                        end
                        else begin
                            $display(";A 2489");		//(= (bv-comp P1_P2_P2_ReadRequest  0b1)   0b0)) ;2489
                            P1_P2_P2_W_R_n <= #1 1'b1; $display(";A 2491");		//(= P1_P2_P2_W_R_n    0b1)) ;2491
                        end
                        if ((P1_P2_P2_CodeFetch == 1'b1)) begin
                            $display(";A 2492");		//(= (bv-comp P1_P2_P2_CodeFetch  0b1)   0b1)) ;2492
                            P1_P2_P2_D_C_n <= #1 1'b0; $display(";A 2494");		//(= P1_P2_P2_D_C_n    0b0)) ;2494
                        end
                        else begin
                            $display(";A 2493");		//(= (bv-comp P1_P2_P2_CodeFetch  0b1)   0b0)) ;2493
                            P1_P2_P2_D_C_n <= #1 1'b1; $display(";A 2495");		//(= P1_P2_P2_D_C_n    0b1)) ;2495
                        end
                        P1_P2_P2_ADS_n <= #1 1'b0; $display(";A 2496");		//(= P1_P2_P2_ADS_n    0b0)) ;2496
                        if ((P1_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 2497");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2497
                            P1_P2_P2_State <= #1 3'sb100; $display(";A 2499");		//(= P1_P2_P2_State    0b100)) ;2499
                        end
                        else begin
                            $display(";A 2498");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2498
                            P1_P2_P2_State <= #1 3'sb110; $display(";A 2500");		//(= P1_P2_P2_State    0b110)) ;2500
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 2501");		//(= P1_P2_P2_State    0b111)) ;2501
                        if ((((P1_P2_P2_READY_n == 1'b1) & (P1_P2_P2_RequestPending == 1'b1)) & (P1_P2_P2_HOLD == 1'b0))) begin
                            $display(";A 2502");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b1) (bv-comp P1_P2_P2_RequestPending  0b1)) (bv-comp P1_P2_P2_HOLD  0b0))   0b1)) ;2502
                            P1_P2_P2_State <= #1 3'sb110; $display(";A 2504");		//(= P1_P2_P2_State    0b110)) ;2504
                        end
                        else begin
                            $display(";A 2503");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b1) (bv-comp P1_P2_P2_RequestPending  0b1)) (bv-comp P1_P2_P2_HOLD  0b0))   0b0)) ;2503
                            if (((P1_P2_P2_READY_n == 1'b0) & (P1_P2_P2_HOLD == 1'b1))) begin
                                $display(";A 2505");		//(= (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b1))   0b1)) ;2505
                                P1_P2_P2_State <= #1 3'sb101; $display(";A 2507");		//(= P1_P2_P2_State    0b101)) ;2507
                            end
                            else begin
                                $display(";A 2506");		//(= (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b1))   0b0)) ;2506
                                if ((((P1_P2_P2_READY_n == 1'b0) & (P1_P2_P2_HOLD == 1'b0)) & (P1_P2_P2_RequestPending == 1'b1))) begin
                                    $display(";A 2508");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b1))   0b1)) ;2508
                                    P1_P2_P2_State <= #1 3'sb010; $display(";A 2510");		//(= P1_P2_P2_State    0b010)) ;2510
                                end
                                else begin
                                    $display(";A 2509");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b1))   0b0)) ;2509
                                    if ((((P1_P2_P2_READY_n == 1'b0) & (P1_P2_P2_HOLD == 1'b0)) & (P1_P2_P2_RequestPending == 1'b0))) begin
                                        $display(";A 2511");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b0))   0b1)) ;2511
                                        P1_P2_P2_State <= #1 3'sb001; $display(";A 2513");		//(= P1_P2_P2_State    0b001)) ;2513
                                    end
                                    else begin
                                        $display(";A 2512");		//(= (bv-and (bv-and (bv-comp P1_P2_P2_READY_n  0b0) (bv-comp P1_P2_P2_HOLD  0b0)) (bv-comp P1_P2_P2_RequestPending  0b0))   0b0)) ;2512
                                        P1_P2_P2_State <= #1 3'sb111; $display(";A 2514");		//(= P1_P2_P2_State    0b111)) ;2514
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:3730
    always @(posedge P1_P2_P2_RESET or posedge P1_P2_P2_CLOCK) begin
        if ((P1_P2_P2_RESET == 1'b1)) begin
            $display(";A 2515");		//(= (bv-comp P1_P2_P2_RESET  0b1)   0b1)) ;2515
            P1_P2_P2_State2 = 4'sb0000; $display(";A 2517");		//(= P1_P2_P2_State2    0b0000)) ;2517
            P1_P2_P2_InstQueue[0] = 8'b00000000; $display(";A 2518");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2518
            P1_P2_P2_InstQueue[1] = 8'b00000000; $display(";A 2519");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2519
            P1_P2_P2_InstQueue[2] = 8'b00000000; $display(";A 2520");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2520
            P1_P2_P2_InstQueue[3] = 8'b00000000; $display(";A 2521");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2521
            P1_P2_P2_InstQueue[4] = 8'b00000000; $display(";A 2522");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2522
            P1_P2_P2_InstQueue[5] = 8'b00000000; $display(";A 2523");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2523
            P1_P2_P2_InstQueue[6] = 8'b00000000; $display(";A 2524");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2524
            P1_P2_P2_InstQueue[7] = 8'b00000000; $display(";A 2525");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2525
            P1_P2_P2_InstQueue[8] = 8'b00000000; $display(";A 2526");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2526
            P1_P2_P2_InstQueue[9] = 8'b00000000; $display(";A 2527");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2527
            P1_P2_P2_InstQueue[10] = 8'b00000000; $display(";A 2528");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2528
            P1_P2_P2_InstQueue[11] = 8'b00000000; $display(";A 2529");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2529
            P1_P2_P2_InstQueue[12] = 8'b00000000; $display(";A 2530");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2530
            P1_P2_P2_InstQueue[13] = 8'b00000000; $display(";A 2531");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2531
            P1_P2_P2_InstQueue[14] = 8'b00000000; $display(";A 2532");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2532
            P1_P2_P2_InstQueue[15] = 8'b00000000; $display(";A 2533");		//(= P1_P2_P2_InstQueue    0b00000000)) ;2533
            P1_P2_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 2534");		//(= P1_P2_P2_InstQueueRd_Addr    0b00000)) ;2534
            P1_P2_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 2535");		//(= P1_P2_P2_InstQueueWr_Addr    0b00000)) ;2535
            P1_P2_P2_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 2536");		//(= P1_P2_P2_InstAddrPointer    0b00000000000000000000000000000000)) ;2536
            P1_P2_P2_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 2537");		//(= P1_P2_P2_PhyAddrPointer    0b00000000000000000000000000000000)) ;2537
            P1_P2_P2_Extended = 1'b0; $display(";A 2538");		//(= P1_P2_P2_Extended    0b0)) ;2538
            P1_P2_P2_More = 1'b0; $display(";A 2539");		//(= P1_P2_P2_More    0b0)) ;2539
            P1_P2_P2_Flush = 1'b0; $display(";A 2540");		//(= P1_P2_P2_Flush    0b0)) ;2540
            P1_P2_P2_lWord = 16'sb0000000000000000; $display(";A 2541");		//(= P1_P2_P2_lWord    0b0000000000000000)) ;2541
            P1_P2_P2_uWord = 15'sb000000000000000; $display(";A 2542");		//(= P1_P2_P2_uWord    0b000000000000000)) ;2542
            P1_P2_P2_fWord = 32'sb00000000000000000000000000000000; $display(";A 2543");		//(= P1_P2_P2_fWord    0b00000000000000000000000000000000)) ;2543
            P1_P2_P2_CodeFetch <= #1 1'b0; $display(";A 2544");		//(= P1_P2_P2_CodeFetch    0b0)) ;2544
            P1_P2_P2_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 2545");		//(= P1_P2_P2_Datao    0b00000000000000000000000000000000)) ;2545
            P1_P2_P2_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 2546");		//(= P1_P2_P2_EAX    0b00000000000000000000000000000000)) ;2546
            P1_P2_P2_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 2547");		//(= P1_P2_P2_EBX    0b00000000000000000000000000000000)) ;2547
            P1_P2_P2_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 2548");		//(= P1_P2_P2_rEIP    0b00000000000000000000000000000000)) ;2548
            P1_P2_P2_ReadRequest <= #1 1'b0; $display(";A 2549");		//(= P1_P2_P2_ReadRequest    0b0)) ;2549
            P1_P2_P2_MemoryFetch <= #1 1'b0; $display(";A 2550");		//(= P1_P2_P2_MemoryFetch    0b0)) ;2550
            P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2551");		//(= P1_P2_P2_RequestPending    0b0)) ;2551
        end
        else begin
            $display(";A 2516");		//(= (bv-comp P1_P2_P2_RESET  0b1)   0b0)) ;2516
            case (P1_P2_P2_State2)
                4'b0000 :
                    begin
                        $display(";A 2552");		//(= P1_P2_P2_State2    0b0000)) ;2552
                        P1_P2_P2_PhyAddrPointer = P1_P2_P2_rEIP; $display(";A 2553");		//(= P1_P2_P2_PhyAddrPointer    P1_P2_P2_rEIP )) ;2553
                        P1_P2_P2_InstAddrPointer = P1_P2_P2_PhyAddrPointer; $display(";A 2554");		//(= P1_P2_P2_InstAddrPointer    P1_P2_P2_PhyAddrPointer )) ;2554
                        P1_P2_P2_State2 = 4'sb0001; $display(";A 2555");		//(= P1_P2_P2_State2    0b0001)) ;2555
                        P1_P2_P2_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 2556");		//(= P1_P2_P2_rEIP    0b00000000000011111111111111110000)) ;2556
                        P1_P2_P2_ReadRequest <= #1 1'b1; $display(";A 2557");		//(= P1_P2_P2_ReadRequest    0b1)) ;2557
                        P1_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 2558");		//(= P1_P2_P2_MemoryFetch    0b1)) ;2558
                        P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2559");		//(= P1_P2_P2_RequestPending    0b1)) ;2559
                    end
                4'b0001 :
                    begin
                        $display(";A 2560");		//(= P1_P2_P2_State2    0b0001)) ;2560
                        P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2561");		//(= P1_P2_P2_RequestPending    0b1)) ;2561
                        P1_P2_P2_ReadRequest <= #1 1'b1; $display(";A 2562");		//(= P1_P2_P2_ReadRequest    0b1)) ;2562
                        P1_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 2563");		//(= P1_P2_P2_MemoryFetch    0b1)) ;2563
                        P1_P2_P2_CodeFetch <= #1 1'b1; $display(";A 2564");		//(= P1_P2_P2_CodeFetch    0b1)) ;2564
                        if ((P1_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 2565");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2565
                            P1_P2_P2_State2 = 4'sb0010; $display(";A 2567");		//(= P1_P2_P2_State2    0b0010)) ;2567
                        end
                        else begin
                            $display(";A 2566");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2566
                            P1_P2_P2_State2 = 4'sb0001; $display(";A 2568");		//(= P1_P2_P2_State2    0b0001)) ;2568
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 2569");		//(= P1_P2_P2_State2    0b0010)) ;2569
                        P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2570");		//(= P1_P2_P2_RequestPending    0b0)) ;2570
                        P1_P2_P2_InstQueue[P1_P2_P2_InstQueueWr_Addr] = (P1_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 2571");		//(= P1_P2_P2_InstQueue    (bv-smod P1_P2_P2_Datai  0b00000000000000000000000100000000))) ;2571
                        P1_P2_P2_InstQueueWr_Addr = ((P1_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2572");		//(= P1_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2572
                        P1_P2_P2_InstQueue[P1_P2_P2_InstQueueWr_Addr] = (P1_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 2573");		//(= P1_P2_P2_InstQueue    (bv-smod P1_P2_P2_Datai  0b00000000000000000000000100000000))) ;2573
                        P1_P2_P2_InstQueueWr_Addr = ((P1_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2574");		//(= P1_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2574
                        if ((P1_P2_P2_StateBS16 == 1'b1)) begin
                            $display(";A 2575");		//(= (bv-comp P1_P2_P2_StateBS16  0b1)   0b1)) ;2575
                            P1_P2_P2_InstQueue[P1_P2_P2_InstQueueWr_Addr] = ((P1_P2_P2_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 2577");		//(= P1_P2_P2_InstQueue    (bv-smod (bv-sdiv P1_P2_P2_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;2577
                            P1_P2_P2_InstQueueWr_Addr = ((P1_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2578");		//(= P1_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2578
                            P1_P2_P2_InstQueue[P1_P2_P2_InstQueueWr_Addr] = ((P1_P2_P2_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 2579");		//(= P1_P2_P2_InstQueue    (bv-smod (bv-sdiv P1_P2_P2_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;2579
                            P1_P2_P2_InstQueueWr_Addr = ((P1_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2580");		//(= P1_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2580
                            P1_P2_P2_PhyAddrPointer = (P1_P2_P2_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 2581");		//(= P1_P2_P2_PhyAddrPointer    (bv-add P1_P2_P2_PhyAddrPointer  0b00000000000000000000000000000100))) ;2581
                            P1_P2_P2_State2 = 4'sb0101; $display(";A 2582");		//(= P1_P2_P2_State2    0b0101)) ;2582
                        end
                        else begin
                            $display(";A 2576");		//(= (bv-comp P1_P2_P2_StateBS16  0b1)   0b0)) ;2576
                            P1_P2_P2_PhyAddrPointer = (P1_P2_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2583");		//(= P1_P2_P2_PhyAddrPointer    (bv-add P1_P2_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;2583
                            if ((P1_P2_P2_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 2584");		//(= (bool-to-bv (bv-slt P1_P2_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;2584
                                P1_P2_P2_rEIP <= #1 (-P1_P2_P2_PhyAddrPointer); $display(";A 2586");		//(= P1_P2_P2_rEIP    (bv-neg P1_P2_P2_PhyAddrPointer ))) ;2586
                            end
                            else begin
                                $display(";A 2585");		//(= (bool-to-bv (bv-slt P1_P2_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;2585
                                P1_P2_P2_rEIP <= #1 P1_P2_P2_PhyAddrPointer; $display(";A 2587");		//(= P1_P2_P2_rEIP    P1_P2_P2_PhyAddrPointer )) ;2587
                            end
                            P1_P2_P2_State2 = 4'sb0011; $display(";A 2588");		//(= P1_P2_P2_State2    0b0011)) ;2588
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 2589");		//(= P1_P2_P2_State2    0b0011)) ;2589
                        P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2590");		//(= P1_P2_P2_RequestPending    0b1)) ;2590
                        if ((P1_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 2591");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2591
                            P1_P2_P2_State2 = 4'sb0100; $display(";A 2593");		//(= P1_P2_P2_State2    0b0100)) ;2593
                        end
                        else begin
                            $display(";A 2592");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2592
                            P1_P2_P2_State2 = 4'sb0011; $display(";A 2594");		//(= P1_P2_P2_State2    0b0011)) ;2594
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 2595");		//(= P1_P2_P2_State2    0b0100)) ;2595
                        P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2596");		//(= P1_P2_P2_RequestPending    0b0)) ;2596
                        P1_P2_P2_InstQueue[P1_P2_P2_InstQueueWr_Addr] = (P1_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 2597");		//(= P1_P2_P2_InstQueue    (bv-smod P1_P2_P2_Datai  0b00000000000000000000000100000000))) ;2597
                        P1_P2_P2_InstQueueWr_Addr = ((P1_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2598");		//(= P1_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2598
                        P1_P2_P2_InstQueue[P1_P2_P2_InstQueueWr_Addr] = (P1_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 2599");		//(= P1_P2_P2_InstQueue    (bv-smod P1_P2_P2_Datai  0b00000000000000000000000100000000))) ;2599
                        P1_P2_P2_InstQueueWr_Addr = ((P1_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2600");		//(= P1_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2600
                        P1_P2_P2_PhyAddrPointer = (P1_P2_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2601");		//(= P1_P2_P2_PhyAddrPointer    (bv-add P1_P2_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;2601
                        P1_P2_P2_State2 = 4'sb0101; $display(";A 2602");		//(= P1_P2_P2_State2    0b0101)) ;2602
                    end
                4'b0101 :
                    begin
                        $display(";A 2603");		//(= P1_P2_P2_State2    0b0101)) ;2603
                        case (P1_P2_P2_InstQueue[P1_P2_P2_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 2604");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b10010000)) ;2604
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2605");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2605
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2606");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2606
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2607");		//(= P1_P2_P2_Flush    0b0)) ;2607
                                    P1_P2_P2_More = 1'b0; $display(";A 2608");		//(= P1_P2_P2_More    0b0)) ;2608
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 2609");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b01100110)) ;2609
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2610");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2610
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2611");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2611
                                    P1_P2_P2_Extended = 1'b1; $display(";A 2612");		//(= P1_P2_P2_Extended    0b1)) ;2612
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2613");		//(= P1_P2_P2_Flush    0b0)) ;2613
                                    P1_P2_P2_More = 1'b0; $display(";A 2614");		//(= P1_P2_P2_More    0b0)) ;2614
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 2615");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b11101011)) ;2615
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 2616");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;2616
                                        if ((P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 2618");		//(= (bool-to-bv (bv-gt P1_P2_P2_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;2618
                                            P1_P2_P2_PhyAddrPointer = ((P1_P2_P2_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 2620");		//(= P1_P2_P2_PhyAddrPointer    (bv-sub (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P1_P2_P2_InstQueue 0 )))) ;2620
                                            P1_P2_P2_InstAddrPointer = P1_P2_P2_PhyAddrPointer; $display(";A 2621");		//(= P1_P2_P2_InstAddrPointer    P1_P2_P2_PhyAddrPointer )) ;2621
                                        end
                                        else begin
                                            $display(";A 2619");		//(= (bool-to-bv (bv-gt P1_P2_P2_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;2619
                                            P1_P2_P2_PhyAddrPointer = ((P1_P2_P2_InstAddrPointer + 32'b00000000000000000000000000000010) + P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 2622");		//(= P1_P2_P2_PhyAddrPointer    (bv-add (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000010) P1_P2_P2_InstQueue 0 ))) ;2622
                                            P1_P2_P2_InstAddrPointer = P1_P2_P2_PhyAddrPointer; $display(";A 2623");		//(= P1_P2_P2_InstAddrPointer    P1_P2_P2_PhyAddrPointer )) ;2623
                                        end
                                        P1_P2_P2_Flush = 1'b1; $display(";A 2624");		//(= P1_P2_P2_Flush    0b1)) ;2624
                                        P1_P2_P2_More = 1'b0; $display(";A 2625");		//(= P1_P2_P2_More    0b0)) ;2625
                                    end
                                    else begin
                                        $display(";A 2617");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;2617
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2626");		//(= P1_P2_P2_Flush    0b0)) ;2626
                                        P1_P2_P2_More = 1'b1; $display(";A 2627");		//(= P1_P2_P2_More    0b1)) ;2627
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 2628");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b11101001)) ;2628
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 2629");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;2629
                                        P1_P2_P2_PhyAddrPointer = ((P1_P2_P2_InstAddrPointer + 32'b00000000000000000000000000000101) + P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 2631");		//(= P1_P2_P2_PhyAddrPointer    (bv-add (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000101) P1_P2_P2_InstQueue 0 ))) ;2631
                                        P1_P2_P2_InstAddrPointer = P1_P2_P2_PhyAddrPointer; $display(";A 2632");		//(= P1_P2_P2_InstAddrPointer    P1_P2_P2_PhyAddrPointer )) ;2632
                                        P1_P2_P2_Flush = 1'b1; $display(";A 2633");		//(= P1_P2_P2_Flush    0b1)) ;2633
                                        P1_P2_P2_More = 1'b0; $display(";A 2634");		//(= P1_P2_P2_More    0b0)) ;2634
                                    end
                                    else begin
                                        $display(";A 2630");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;2630
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2635");		//(= P1_P2_P2_Flush    0b0)) ;2635
                                        P1_P2_P2_More = 1'b1; $display(";A 2636");		//(= P1_P2_P2_More    0b1)) ;2636
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 2637");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b11101010)) ;2637
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2638");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2638
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2639");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2639
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2640");		//(= P1_P2_P2_Flush    0b0)) ;2640
                                    P1_P2_P2_More = 1'b0; $display(";A 2641");		//(= P1_P2_P2_More    0b0)) ;2641
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 2642");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b10110000)) ;2642
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2643");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2643
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2644");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2644
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2645");		//(= P1_P2_P2_Flush    0b0)) ;2645
                                    P1_P2_P2_More = 1'b0; $display(";A 2646");		//(= P1_P2_P2_More    0b0)) ;2646
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 2647");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b10111000)) ;2647
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 2648");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;2648
                                        P1_P2_P2_EAX <= #1 ((((P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 2650");		//(= P1_P2_P2_EAX    (bv-add (bv-add (bv-add (bv-mul P1_P2_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P2_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P2_P2_InstQueue 0  0b00000000000000000000000100000000)) P1_P2_P2_InstQueue 0 ))) ;2650
                                        P1_P2_P2_More = 1'b0; $display(";A 2651");		//(= P1_P2_P2_More    0b0)) ;2651
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2652");		//(= P1_P2_P2_Flush    0b0)) ;2652
                                        P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 2653");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;2653
                                        P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 2654");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;2654
                                    end
                                    else begin
                                        $display(";A 2649");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;2649
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2655");		//(= P1_P2_P2_Flush    0b0)) ;2655
                                        P1_P2_P2_More = 1'b1; $display(";A 2656");		//(= P1_P2_P2_More    0b1)) ;2656
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 2657");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b10111011)) ;2657
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 2658");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;2658
                                        P1_P2_P2_EBX <= #1 ((((P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P2_P2_InstQueue[((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 2660");		//(= P1_P2_P2_EBX    (bv-add (bv-add (bv-add (bv-mul P1_P2_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P2_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P2_P2_InstQueue 0  0b00000000000000000000000100000000)) P1_P2_P2_InstQueue 0 ))) ;2660
                                        P1_P2_P2_More = 1'b0; $display(";A 2661");		//(= P1_P2_P2_More    0b0)) ;2661
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2662");		//(= P1_P2_P2_Flush    0b0)) ;2662
                                        P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 2663");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;2663
                                        P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 2664");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;2664
                                    end
                                    else begin
                                        $display(";A 2659");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;2659
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2665");		//(= P1_P2_P2_Flush    0b0)) ;2665
                                        P1_P2_P2_More = 1'b1; $display(";A 2666");		//(= P1_P2_P2_More    0b1)) ;2666
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 2667");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b10001011)) ;2667
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2668");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2668
                                        if ((P1_P2_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 2670");		//(= (bool-to-bv (bv-slt P1_P2_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;2670
                                            P1_P2_P2_rEIP <= #1 (-P1_P2_P2_EBX); $display(";A 2672");		//(= P1_P2_P2_rEIP    (bv-neg P1_P2_P2_EBX ))) ;2672
                                        end
                                        else begin
                                            $display(";A 2671");		//(= (bool-to-bv (bv-slt P1_P2_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;2671
                                            P1_P2_P2_rEIP <= #1 P1_P2_P2_EBX; $display(";A 2673");		//(= P1_P2_P2_rEIP    P1_P2_P2_EBX )) ;2673
                                        end
                                        P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2674");		//(= P1_P2_P2_RequestPending    0b1)) ;2674
                                        P1_P2_P2_ReadRequest <= #1 1'b1; $display(";A 2675");		//(= P1_P2_P2_ReadRequest    0b1)) ;2675
                                        P1_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 2676");		//(= P1_P2_P2_MemoryFetch    0b1)) ;2676
                                        P1_P2_P2_CodeFetch <= #1 1'b0; $display(";A 2677");		//(= P1_P2_P2_CodeFetch    0b0)) ;2677
                                        if ((P1_P2_P2_READY_n == 1'b0)) begin
                                            $display(";A 2678");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2678
                                            P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2680");		//(= P1_P2_P2_RequestPending    0b0)) ;2680
                                            P1_P2_P2_uWord = (P1_P2_P2_Datai % 32'b00000000000000001000000000000000); $display(";A 2681");		//(= P1_P2_P2_uWord    (bv-smod P1_P2_P2_Datai  0b00000000000000001000000000000000))) ;2681
                                            if ((P1_P2_P2_StateBS16 == 1'b1)) begin
                                                $display(";A 2682");		//(= (bv-comp P1_P2_P2_StateBS16  0b1)   0b1)) ;2682
                                                P1_P2_P2_lWord = (P1_P2_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 2684");		//(= P1_P2_P2_lWord    (bv-smod P1_P2_P2_Datai  0b00000000000000010000000000000000))) ;2684
                                            end
                                            else begin
                                                $display(";A 2683");		//(= (bv-comp P1_P2_P2_StateBS16  0b1)   0b0)) ;2683
                                                P1_P2_P2_rEIP <= #1 (P1_P2_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 2685");		//(= P1_P2_P2_rEIP    (bv-add P1_P2_P2_rEIP  0b00000000000000000000000000000010))) ;2685
                                                P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2686");		//(= P1_P2_P2_RequestPending    0b1)) ;2686
                                                if ((P1_P2_P2_READY_n == 1'b0)) begin
                                                    $display(";A 2687");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2687
                                                    P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2689");		//(= P1_P2_P2_RequestPending    0b0)) ;2689
                                                    P1_P2_P2_lWord = (P1_P2_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 2690");		//(= P1_P2_P2_lWord    (bv-smod P1_P2_P2_Datai  0b00000000000000010000000000000000))) ;2690
                                                end
                                                else begin
                                                    $display(";A 2688");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2688
                                                end
                                            end
                                            if ((P1_P2_P2_READY_n == 1'b0)) begin
                                                $display(";A 2691");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2691
                                                P1_P2_P2_EAX <= #1 ((P1_P2_P2_uWord * 32'b00000000000000010000000000000000) + P1_P2_P2_lWord); $display(";A 2693");		//(= P1_P2_P2_EAX    (bv-add (bv-mul P1_P2_P2_uWord  0b00000000000000010000000000000000) P1_P2_P2_lWord ))) ;2693
                                                P1_P2_P2_More = 1'b0; $display(";A 2694");		//(= P1_P2_P2_More    0b0)) ;2694
                                                P1_P2_P2_Flush = 1'b0; $display(";A 2695");		//(= P1_P2_P2_Flush    0b0)) ;2695
                                                P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2696");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;2696
                                                P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2697");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2697
                                            end
                                            else begin
                                                $display(";A 2692");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2692
                                            end
                                        end
                                        else begin
                                            $display(";A 2679");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2679
                                        end
                                    end
                                    else begin
                                        $display(";A 2669");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2669
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2698");		//(= P1_P2_P2_Flush    0b0)) ;2698
                                        P1_P2_P2_More = 1'b1; $display(";A 2699");		//(= P1_P2_P2_More    0b1)) ;2699
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 2700");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b10001001)) ;2700
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2701");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2701
                                        if ((P1_P2_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 2703");		//(= (bool-to-bv (bv-slt P1_P2_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;2703
                                            P1_P2_P2_rEIP <= #1 P1_P2_P2_EBX; $display(";A 2705");		//(= P1_P2_P2_rEIP    P1_P2_P2_EBX )) ;2705
                                        end
                                        else begin
                                            $display(";A 2704");		//(= (bool-to-bv (bv-slt P1_P2_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;2704
                                            P1_P2_P2_rEIP <= #1 P1_P2_P2_EBX; $display(";A 2706");		//(= P1_P2_P2_rEIP    P1_P2_P2_EBX )) ;2706
                                        end
                                        P1_P2_P2_lWord = (P1_P2_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 2707");		//(= P1_P2_P2_lWord    (bv-smod P1_P2_P2_EAX  0b00000000000000010000000000000000))) ;2707
                                        P1_P2_P2_uWord = ((P1_P2_P2_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 2708");		//(= P1_P2_P2_uWord    (bv-smod (bv-sdiv P1_P2_P2_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;2708
                                        P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2709");		//(= P1_P2_P2_RequestPending    0b1)) ;2709
                                        P1_P2_P2_ReadRequest <= #1 1'b0; $display(";A 2710");		//(= P1_P2_P2_ReadRequest    0b0)) ;2710
                                        P1_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 2711");		//(= P1_P2_P2_MemoryFetch    0b1)) ;2711
                                        P1_P2_P2_CodeFetch <= #1 1'b0; $display(";A 2712");		//(= P1_P2_P2_CodeFetch    0b0)) ;2712
                                        if (((P1_P2_P2_State == 32'b00000000000000000000000000000010) | (P1_P2_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 2713");		//(= (bv-or (bv-comp P1_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P2_State  0b00000000000000000000000000000100))   0b1)) ;2713
                                            P1_P2_P2_Datao <= #1 ((P1_P2_P2_uWord * 32'b00000000000000010000000000000000) + P1_P2_P2_lWord); $display(";A 2715");		//(= P1_P2_P2_Datao    (bv-add (bv-mul P1_P2_P2_uWord  0b00000000000000010000000000000000) P1_P2_P2_lWord ))) ;2715
                                            if ((P1_P2_P2_READY_n == 1'b0)) begin
                                                $display(";A 2716");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2716
                                                P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2718");		//(= P1_P2_P2_RequestPending    0b0)) ;2718
                                                if ((P1_P2_P2_StateBS16 == 1'b0)) begin
                                                    $display(";A 2719");		//(= (bv-comp P1_P2_P2_StateBS16  0b0)   0b1)) ;2719
                                                    P1_P2_P2_rEIP <= #1 (P1_P2_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 2721");		//(= P1_P2_P2_rEIP    (bv-add P1_P2_P2_rEIP  0b00000000000000000000000000000010))) ;2721
                                                    P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2722");		//(= P1_P2_P2_RequestPending    0b1)) ;2722
                                                    P1_P2_P2_ReadRequest <= #1 1'b0; $display(";A 2723");		//(= P1_P2_P2_ReadRequest    0b0)) ;2723
                                                    P1_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 2724");		//(= P1_P2_P2_MemoryFetch    0b1)) ;2724
                                                    P1_P2_P2_CodeFetch <= #1 1'b0; $display(";A 2725");		//(= P1_P2_P2_CodeFetch    0b0)) ;2725
                                                    P1_P2_P2_State2 = 4'sb0110; $display(";A 2726");		//(= P1_P2_P2_State2    0b0110)) ;2726
                                                end
                                                else begin
                                                    $display(";A 2720");		//(= (bv-comp P1_P2_P2_StateBS16  0b0)   0b0)) ;2720
                                                end
                                                P1_P2_P2_More = 1'b0; $display(";A 2727");		//(= P1_P2_P2_More    0b0)) ;2727
                                                P1_P2_P2_Flush = 1'b0; $display(";A 2728");		//(= P1_P2_P2_Flush    0b0)) ;2728
                                                P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2729");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;2729
                                                P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2730");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2730
                                            end
                                            else begin
                                                $display(";A 2717");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2717
                                            end
                                        end
                                        else begin
                                            $display(";A 2714");		//(= (bv-or (bv-comp P1_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P2_State  0b00000000000000000000000000000100))   0b0)) ;2714
                                        end
                                    end
                                    else begin
                                        $display(";A 2702");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2702
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2731");		//(= P1_P2_P2_Flush    0b0)) ;2731
                                        P1_P2_P2_More = 1'b1; $display(";A 2732");		//(= P1_P2_P2_More    0b1)) ;2732
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 2733");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b11100100)) ;2733
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2734");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2734
                                        P1_P2_P2_rEIP <= #1 (P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 2736");		//(= P1_P2_P2_rEIP    (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;2736
                                        P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2737");		//(= P1_P2_P2_RequestPending    0b1)) ;2737
                                        P1_P2_P2_ReadRequest <= #1 1'b1; $display(";A 2738");		//(= P1_P2_P2_ReadRequest    0b1)) ;2738
                                        P1_P2_P2_MemoryFetch <= #1 1'b0; $display(";A 2739");		//(= P1_P2_P2_MemoryFetch    0b0)) ;2739
                                        P1_P2_P2_CodeFetch <= #1 1'b0; $display(";A 2740");		//(= P1_P2_P2_CodeFetch    0b0)) ;2740
                                        if ((P1_P2_P2_READY_n == 1'b0)) begin
                                            $display(";A 2741");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2741
                                            P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2743");		//(= P1_P2_P2_RequestPending    0b0)) ;2743
                                            P1_P2_P2_EAX <= #1 P1_P2_P2_Datai; $display(";A 2744");		//(= P1_P2_P2_EAX    P1_P2_P2_Datai )) ;2744
                                            P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2745");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;2745
                                            P1_P2_P2_InstQueueRd_Addr = (P1_P2_P2_InstQueueRd_Addr + 5'b00010); $display(";A 2746");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-add P1_P2_P2_InstQueueRd_Addr  0b00010))) ;2746
                                            P1_P2_P2_Flush = 1'b0; $display(";A 2747");		//(= P1_P2_P2_Flush    0b0)) ;2747
                                            P1_P2_P2_More = 1'b0; $display(";A 2748");		//(= P1_P2_P2_More    0b0)) ;2748
                                        end
                                        else begin
                                            $display(";A 2742");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2742
                                        end
                                    end
                                    else begin
                                        $display(";A 2735");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2735
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2749");		//(= P1_P2_P2_Flush    0b0)) ;2749
                                        P1_P2_P2_More = 1'b1; $display(";A 2750");		//(= P1_P2_P2_More    0b1)) ;2750
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 2751");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b11100110)) ;2751
                                    if (((P1_P2_P2_InstQueueWr_Addr - P1_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 2752");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;2752
                                        P1_P2_P2_rEIP <= #1 (P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 2754");		//(= P1_P2_P2_rEIP    (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;2754
                                        P1_P2_P2_RequestPending <= #1 1'b1; $display(";A 2755");		//(= P1_P2_P2_RequestPending    0b1)) ;2755
                                        P1_P2_P2_ReadRequest <= #1 1'b0; $display(";A 2756");		//(= P1_P2_P2_ReadRequest    0b0)) ;2756
                                        P1_P2_P2_MemoryFetch <= #1 1'b0; $display(";A 2757");		//(= P1_P2_P2_MemoryFetch    0b0)) ;2757
                                        P1_P2_P2_CodeFetch <= #1 1'b0; $display(";A 2758");		//(= P1_P2_P2_CodeFetch    0b0)) ;2758
                                        if (((P1_P2_P2_State == 32'b00000000000000000000000000000010) | (P1_P2_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 2759");		//(= (bv-or (bv-comp P1_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P2_State  0b00000000000000000000000000000100))   0b1)) ;2759
                                            P1_P2_P2_fWord = (P1_P2_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 2761");		//(= P1_P2_P2_fWord    (bv-smod P1_P2_P2_EAX  0b00000000000000010000000000000000))) ;2761
                                            P1_P2_P2_Datao <= #1 P1_P2_P2_fWord; $display(";A 2762");		//(= P1_P2_P2_Datao    P1_P2_P2_fWord )) ;2762
                                            if ((P1_P2_P2_READY_n == 1'b0)) begin
                                                $display(";A 2763");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2763
                                                P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2765");		//(= P1_P2_P2_RequestPending    0b0)) ;2765
                                                P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2766");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;2766
                                                P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2767");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2767
                                                P1_P2_P2_Flush = 1'b0; $display(";A 2768");		//(= P1_P2_P2_Flush    0b0)) ;2768
                                                P1_P2_P2_More = 1'b0; $display(";A 2769");		//(= P1_P2_P2_More    0b0)) ;2769
                                            end
                                            else begin
                                                $display(";A 2764");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2764
                                            end
                                        end
                                        else begin
                                            $display(";A 2760");		//(= (bv-or (bv-comp P1_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P2_State  0b00000000000000000000000000000100))   0b0)) ;2760
                                        end
                                    end
                                    else begin
                                        $display(";A 2753");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P2_InstQueueWr_Addr  P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;2753
                                        P1_P2_P2_Flush = 1'b0; $display(";A 2770");		//(= P1_P2_P2_Flush    0b0)) ;2770
                                        P1_P2_P2_More = 1'b1; $display(";A 2771");		//(= P1_P2_P2_More    0b1)) ;2771
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 2772");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b00000100)) ;2772
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2773");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2773
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2774");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2774
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2775");		//(= P1_P2_P2_Flush    0b0)) ;2775
                                    P1_P2_P2_More = 1'b0; $display(";A 2776");		//(= P1_P2_P2_More    0b0)) ;2776
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 2777");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b00000101)) ;2777
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2778");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2778
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2779");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2779
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2780");		//(= P1_P2_P2_Flush    0b0)) ;2780
                                    P1_P2_P2_More = 1'b0; $display(";A 2781");		//(= P1_P2_P2_More    0b0)) ;2781
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 2782");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b11010000)) ;2782
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2783");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;2783
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2784");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2784
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2785");		//(= P1_P2_P2_Flush    0b0)) ;2785
                                    P1_P2_P2_More = 1'b0; $display(";A 2786");		//(= P1_P2_P2_More    0b0)) ;2786
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 2787");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b11000000)) ;2787
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 2788");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;2788
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 2789");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;2789
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2790");		//(= P1_P2_P2_Flush    0b0)) ;2790
                                    P1_P2_P2_More = 1'b0; $display(";A 2791");		//(= P1_P2_P2_More    0b0)) ;2791
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 2792");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b01000000)) ;2792
                                    P1_P2_P2_EAX <= #1 (P1_P2_P2_EAX + 32'sb00000000000000000000000000000001); $display(";A 2793");		//(= P1_P2_P2_EAX    (bv-add P1_P2_P2_EAX  0b00000000000000000000000000000001))) ;2793
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2794");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2794
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2795");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2795
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2796");		//(= P1_P2_P2_Flush    0b0)) ;2796
                                    P1_P2_P2_More = 1'b0; $display(";A 2797");		//(= P1_P2_P2_More    0b0)) ;2797
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 2798");		//(= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr )   0b01000011)) ;2798
                                    P1_P2_P2_EBX <= #1 (P1_P2_P2_EBX + 32'sb00000000000000000000000000000001); $display(";A 2799");		//(= P1_P2_P2_EBX    (bv-add P1_P2_P2_EBX  0b00000000000000000000000000000001))) ;2799
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2800");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2800
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2801");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2801
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2802");		//(= P1_P2_P2_Flush    0b0)) ;2802
                                    P1_P2_P2_More = 1'b0; $display(";A 2803");		//(= P1_P2_P2_More    0b0)) ;2803
                                end
                            default:
                                begin
                                    $display(";A 2804");		//(= (and (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b10010000) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b01100110) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b11101011) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b11101001) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b11101010) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b10110000) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b10111000) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b10111011) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b10001011) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b10001001) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b11100100) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b11100110) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b00000100) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b00000101) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b11010000) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b11000000) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b01000000) (/= ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ) 0b01000011))   true)) ;2804
                                    P1_P2_P2_InstAddrPointer = (P1_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 2805");		//(= P1_P2_P2_InstAddrPointer    (bv-add P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;2805
                                    P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2806");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2806
                                    P1_P2_P2_Flush = 1'b0; $display(";A 2807");		//(= P1_P2_P2_Flush    0b0)) ;2807
                                    P1_P2_P2_More = 1'b0; $display(";A 2808");		//(= P1_P2_P2_More    0b0)) ;2808
                                end
                        endcase
                        if (((~(P1_P2_P2_InstQueueRd_Addr < P1_P2_P2_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P1_P2_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P1_P2_P2_Flush) | P1_P2_P2_More))) begin
                            $display(";A 2809");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P2_P2_InstQueueRd_Addr  P1_P2_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P2_P2_Flush ) P1_P2_P2_More ))   0b1)) ;2809
                            P1_P2_P2_State2 = 4'sb0111; $display(";A 2811");		//(= P1_P2_P2_State2    0b0111)) ;2811
                        end
                        else begin
                            $display(";A 2810");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P2_P2_InstQueueRd_Addr  P1_P2_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P2_P2_Flush ) P1_P2_P2_More ))   0b0)) ;2810
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 2812");		//(= P1_P2_P2_State2    0b0110)) ;2812
                        P1_P2_P2_Datao <= #1 ((P1_P2_P2_uWord * 32'b00000000000000010000000000000000) + P1_P2_P2_lWord); $display(";A 2813");		//(= P1_P2_P2_Datao    (bv-add (bv-mul P1_P2_P2_uWord  0b00000000000000010000000000000000) P1_P2_P2_lWord ))) ;2813
                        if ((P1_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 2814");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b1)) ;2814
                            P1_P2_P2_RequestPending <= #1 1'b0; $display(";A 2816");		//(= P1_P2_P2_RequestPending    0b0)) ;2816
                            P1_P2_P2_State2 = 4'sb0101; $display(";A 2817");		//(= P1_P2_P2_State2    0b0101)) ;2817
                        end
                        else begin
                            $display(";A 2815");		//(= (bv-comp P1_P2_P2_READY_n  0b0)   0b0)) ;2815
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 2818");		//(= P1_P2_P2_State2    0b0111)) ;2818
                        if (P1_P2_P2_Flush) begin
                            $display(";A 2819");		//(= P1_P2_P2_Flush    0b1)) ;2819
                            P1_P2_P2_InstQueueRd_Addr = 5'sb00001; $display(";A 2821");		//(= P1_P2_P2_InstQueueRd_Addr    0b00001)) ;2821
                            P1_P2_P2_InstQueueWr_Addr = 5'sb00001; $display(";A 2822");		//(= P1_P2_P2_InstQueueWr_Addr    0b00001)) ;2822
                            if ((P1_P2_P2_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 2823");		//(= (bool-to-bv (bv-slt P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;2823
                                P1_P2_P2_fWord = (-P1_P2_P2_InstAddrPointer); $display(";A 2825");		//(= P1_P2_P2_fWord    (bv-neg P1_P2_P2_InstAddrPointer ))) ;2825
                            end
                            else begin
                                $display(";A 2824");		//(= (bool-to-bv (bv-slt P1_P2_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;2824
                                P1_P2_P2_fWord = P1_P2_P2_InstAddrPointer; $display(";A 2826");		//(= P1_P2_P2_fWord    P1_P2_P2_InstAddrPointer )) ;2826
                            end
                            if (((P1_P2_P2_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 2827");		//(= (bv-comp (bv-smod P1_P2_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;2827
                                P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + (P1_P2_P2_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 2829");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  (bv-smod P1_P2_P2_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;2829
                            end
                            else begin
                                $display(";A 2828");		//(= (bv-comp (bv-smod P1_P2_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;2828
                            end
                        end
                        else begin
                            $display(";A 2820");		//(= P1_P2_P2_Flush    0b0)) ;2820
                        end
                        if (((32'b00000000000000000000000000001111 - P1_P2_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 2830");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;2830
                            P1_P2_P2_State2 = 4'sb1000; $display(";A 2832");		//(= P1_P2_P2_State2    0b1000)) ;2832
                            P1_P2_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 2833");		//(= P1_P2_P2_InstQueueWr_Addr    0b00000)) ;2833
                        end
                        else begin
                            $display(";A 2831");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;2831
                            P1_P2_P2_State2 = 4'sb1001; $display(";A 2834");		//(= P1_P2_P2_State2    0b1001)) ;2834
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 2835");		//(= P1_P2_P2_State2    0b1000)) ;2835
                        if ((P1_P2_P2_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 2836");		//(= (bool-to-bv (bv-le P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;2836
                            P1_P2_P2_InstQueue[P1_P2_P2_InstQueueWr_Addr] = P1_P2_P2_InstQueue[P1_P2_P2_InstQueueRd_Addr]; $display(";A 2838");		//(= P1_P2_P2_InstQueue    ( P1_P2_P2_InstQueue P1_P2_P2_InstQueueRd_Addr ))) ;2838
                            P1_P2_P2_InstQueueRd_Addr = ((P1_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2839");		//(= P1_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2839
                            P1_P2_P2_InstQueueWr_Addr = ((P1_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 2840");		//(= P1_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;2840
                            P1_P2_P2_State2 = 4'sb1000; $display(";A 2841");		//(= P1_P2_P2_State2    0b1000)) ;2841
                        end
                        else begin
                            $display(";A 2837");		//(= (bool-to-bv (bv-le P1_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;2837
                            P1_P2_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 2842");		//(= P1_P2_P2_InstQueueRd_Addr    0b00000)) ;2842
                            P1_P2_P2_State2 = 4'sb1001; $display(";A 2843");		//(= P1_P2_P2_State2    0b1001)) ;2843
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 2844");		//(= P1_P2_P2_State2    0b1001)) ;2844
                        P1_P2_P2_rEIP <= #1 P1_P2_P2_PhyAddrPointer; $display(";A 2845");		//(= P1_P2_P2_rEIP    P1_P2_P2_PhyAddrPointer )) ;2845
                        P1_P2_P2_State2 = 4'sb0001; $display(";A 2846");		//(= P1_P2_P2_State2    0b0001)) ;2846
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:4169
    always @(posedge P1_P2_P2_RESET or posedge P1_P2_P2_CLOCK) begin
        if ((P1_P2_P2_RESET == 1'b1)) begin
            $display(";A 2847");		//(= (bv-comp P1_P2_P2_RESET  0b1)   0b1)) ;2847
            P1_P2_P2_ByteEnable <= #1 4'b0000; $display(";A 2849");		//(= P1_P2_P2_ByteEnable    0b0000)) ;2849
            P1_P2_P2_NonAligned <= #1 1'b0; $display(";A 2850");		//(= P1_P2_P2_NonAligned    0b0)) ;2850
        end
        else begin
            $display(";A 2848");		//(= (bv-comp P1_P2_P2_RESET  0b1)   0b0)) ;2848
            case (P1_P2_P2_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 2851");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000000)) ;2851
                        case ((P1_P2_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 2852");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;2852
                                    P1_P2_P2_ByteEnable <= #1 4'b1110; $display(";A 2853");		//(= P1_P2_P2_ByteEnable    0b1110)) ;2853
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 2854");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;2854
                                    P1_P2_P2_ByteEnable <= #1 4'b1101; $display(";A 2855");		//(= P1_P2_P2_ByteEnable    0b1101)) ;2855
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 2856");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;2856
                                    P1_P2_P2_ByteEnable <= #1 4'b1011; $display(";A 2857");		//(= P1_P2_P2_ByteEnable    0b1011)) ;2857
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 2858");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;2858
                                    P1_P2_P2_ByteEnable <= #1 4'b0111; $display(";A 2859");		//(= P1_P2_P2_ByteEnable    0b0111)) ;2859
                                end
                            default:
                                begin
                                    $display(";A 2860");		//(= (and (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;2860
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 2861");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000001)) ;2861
                        case ((P1_P2_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 2862");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;2862
                                    P1_P2_P2_ByteEnable <= #1 4'b1100; $display(";A 2863");		//(= P1_P2_P2_ByteEnable    0b1100)) ;2863
                                    P1_P2_P2_NonAligned <= #1 1'b0; $display(";A 2864");		//(= P1_P2_P2_NonAligned    0b0)) ;2864
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 2865");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;2865
                                    P1_P2_P2_ByteEnable <= #1 4'b1001; $display(";A 2866");		//(= P1_P2_P2_ByteEnable    0b1001)) ;2866
                                    P1_P2_P2_NonAligned <= #1 1'b0; $display(";A 2867");		//(= P1_P2_P2_NonAligned    0b0)) ;2867
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 2868");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;2868
                                    P1_P2_P2_ByteEnable <= #1 4'b0011; $display(";A 2869");		//(= P1_P2_P2_ByteEnable    0b0011)) ;2869
                                    P1_P2_P2_NonAligned <= #1 1'b0; $display(";A 2870");		//(= P1_P2_P2_NonAligned    0b0)) ;2870
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 2871");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;2871
                                    P1_P2_P2_ByteEnable <= #1 4'b0111; $display(";A 2872");		//(= P1_P2_P2_ByteEnable    0b0111)) ;2872
                                    P1_P2_P2_NonAligned <= #1 1'b1; $display(";A 2873");		//(= P1_P2_P2_NonAligned    0b1)) ;2873
                                end
                            default:
                                begin
                                    $display(";A 2874");		//(= (and (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;2874
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 2875");		//(= P1_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;2875
                        case ((P1_P2_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 2876");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;2876
                                    P1_P2_P2_ByteEnable <= #1 4'b0000; $display(";A 2877");		//(= P1_P2_P2_ByteEnable    0b0000)) ;2877
                                    P1_P2_P2_NonAligned <= #1 1'b0; $display(";A 2878");		//(= P1_P2_P2_NonAligned    0b0)) ;2878
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 2879");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;2879
                                    P1_P2_P2_ByteEnable <= #1 4'b0001; $display(";A 2880");		//(= P1_P2_P2_ByteEnable    0b0001)) ;2880
                                    P1_P2_P2_NonAligned <= #1 1'b1; $display(";A 2881");		//(= P1_P2_P2_NonAligned    0b1)) ;2881
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 2882");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;2882
                                    P1_P2_P2_NonAligned <= #1 1'b1; $display(";A 2883");		//(= P1_P2_P2_NonAligned    0b1)) ;2883
                                    P1_P2_P2_ByteEnable <= #1 4'b0011; $display(";A 2884");		//(= P1_P2_P2_ByteEnable    0b0011)) ;2884
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 2885");		//(= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;2885
                                    P1_P2_P2_NonAligned <= #1 1'b1; $display(";A 2886");		//(= P1_P2_P2_NonAligned    0b1)) ;2886
                                    P1_P2_P2_ByteEnable <= #1 4'b0111; $display(";A 2887");		//(= P1_P2_P2_ByteEnable    0b0111)) ;2887
                                end
                            default:
                                begin
                                    $display(";A 2888");		//(= (and (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;2888
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 2889");		//(= (and (/= P1_P2_P2_DataWidth  0b00000000000000000000000000000000) (/= P1_P2_P2_DataWidth  0b00000000000000000000000000000001) (/= P1_P2_P2_DataWidth  0b00000000000000000000000000000010))   true)) ;2889
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:4357
    always @(posedge P1_P2_P3_RESET or posedge P1_P2_P3_CLOCK) begin
        if ((P1_P2_P3_RESET == 1'b1)) begin
            $display(";A 2890");		//(= (bv-comp P1_P2_P3_RESET  0b1)   0b1)) ;2890
            P1_P2_P3_BE_n <= #1 4'b0000; $display(";A 2892");		//(= P1_P2_P3_BE_n    0b0000)) ;2892
            P1_P2_P3_Address <= #1 30'sb000000000000000000000000000000; $display(";A 2893");		//(= P1_P2_P3_Address    0b000000000000000000000000000000)) ;2893
            P1_P2_P3_W_R_n <= #1 1'b0; $display(";A 2894");		//(= P1_P2_P3_W_R_n    0b0)) ;2894
            P1_P2_P3_D_C_n <= #1 1'b0; $display(";A 2895");		//(= P1_P2_P3_D_C_n    0b0)) ;2895
            P1_P2_P3_M_IO_n <= #1 1'b0; $display(";A 2896");		//(= P1_P2_P3_M_IO_n    0b0)) ;2896
            P1_P2_P3_ADS_n <= #1 1'b0; $display(";A 2897");		//(= P1_P2_P3_ADS_n    0b0)) ;2897
            P1_P2_P3_State <= #1 3'sb000; $display(";A 2898");		//(= P1_P2_P3_State    0b000)) ;2898
            P1_P2_P3_StateNA <= #1 1'b0; $display(";A 2899");		//(= P1_P2_P3_StateNA    0b0)) ;2899
            P1_P2_P3_StateBS16 <= #1 1'b0; $display(";A 2900");		//(= P1_P2_P3_StateBS16    0b0)) ;2900
            P1_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 2901");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000000)) ;2901
        end
        else begin
            $display(";A 2891");		//(= (bv-comp P1_P2_P3_RESET  0b1)   0b0)) ;2891
            case (P1_P2_P3_State)
                3'b000 :
                    begin
                        $display(";A 2902");		//(= P1_P2_P3_State    0b000)) ;2902
                        P1_P2_P3_D_C_n <= #1 1'b1; $display(";A 2903");		//(= P1_P2_P3_D_C_n    0b1)) ;2903
                        P1_P2_P3_ADS_n <= #1 1'b1; $display(";A 2904");		//(= P1_P2_P3_ADS_n    0b1)) ;2904
                        P1_P2_P3_State <= #1 3'sb001; $display(";A 2905");		//(= P1_P2_P3_State    0b001)) ;2905
                        P1_P2_P3_StateNA <= #1 1'b1; $display(";A 2906");		//(= P1_P2_P3_StateNA    0b1)) ;2906
                        P1_P2_P3_StateBS16 <= #1 1'b1; $display(";A 2907");		//(= P1_P2_P3_StateBS16    0b1)) ;2907
                        P1_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 2908");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;2908
                        P1_P2_P3_State <= #1 3'sb001; $display(";A 2909");		//(= P1_P2_P3_State    0b001)) ;2909
                    end
                3'b001 :
                    begin
                        $display(";A 2910");		//(= P1_P2_P3_State    0b001)) ;2910
                        if ((P1_P2_P3_RequestPending == 1'b1)) begin
                            $display(";A 2911");		//(= (bv-comp P1_P2_P3_RequestPending  0b1)   0b1)) ;2911
                            P1_P2_P3_State <= #1 3'sb010; $display(";A 2913");		//(= P1_P2_P3_State    0b010)) ;2913
                        end
                        else begin
                            $display(";A 2912");		//(= (bv-comp P1_P2_P3_RequestPending  0b1)   0b0)) ;2912
                            if ((P1_P2_P3_HOLD == 1'b1)) begin
                                $display(";A 2914");		//(= (bv-comp P1_P2_P3_HOLD  0b1)   0b1)) ;2914
                                P1_P2_P3_State <= #1 3'sb101; $display(";A 2916");		//(= P1_P2_P3_State    0b101)) ;2916
                            end
                            else begin
                                $display(";A 2915");		//(= (bv-comp P1_P2_P3_HOLD  0b1)   0b0)) ;2915
                                P1_P2_P3_State <= #1 3'sb001; $display(";A 2917");		//(= P1_P2_P3_State    0b001)) ;2917
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 2918");		//(= P1_P2_P3_State    0b010)) ;2918
                        P1_P2_P3_Address <= #1 ((P1_P2_P3_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 2919");		//(= P1_P2_P3_Address    (bv-smod (bv-sdiv P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;2919
                        P1_P2_P3_BE_n <= #1 P1_P2_P3_ByteEnable; $display(";A 2920");		//(= P1_P2_P3_BE_n    P1_P2_P3_ByteEnable )) ;2920
                        P1_P2_P3_M_IO_n <= #1 P1_P2_P3_MemoryFetch; $display(";A 2921");		//(= P1_P2_P3_M_IO_n    P1_P2_P3_MemoryFetch )) ;2921
                        if ((P1_P2_P3_ReadRequest == 1'b1)) begin
                            $display(";A 2922");		//(= (bv-comp P1_P2_P3_ReadRequest  0b1)   0b1)) ;2922
                            P1_P2_P3_W_R_n <= #1 1'b0; $display(";A 2924");		//(= P1_P2_P3_W_R_n    0b0)) ;2924
                        end
                        else begin
                            $display(";A 2923");		//(= (bv-comp P1_P2_P3_ReadRequest  0b1)   0b0)) ;2923
                            P1_P2_P3_W_R_n <= #1 1'b1; $display(";A 2925");		//(= P1_P2_P3_W_R_n    0b1)) ;2925
                        end
                        if ((P1_P2_P3_CodeFetch == 1'b1)) begin
                            $display(";A 2926");		//(= (bv-comp P1_P2_P3_CodeFetch  0b1)   0b1)) ;2926
                            P1_P2_P3_D_C_n <= #1 1'b0; $display(";A 2928");		//(= P1_P2_P3_D_C_n    0b0)) ;2928
                        end
                        else begin
                            $display(";A 2927");		//(= (bv-comp P1_P2_P3_CodeFetch  0b1)   0b0)) ;2927
                            P1_P2_P3_D_C_n <= #1 1'b1; $display(";A 2929");		//(= P1_P2_P3_D_C_n    0b1)) ;2929
                        end
                        P1_P2_P3_ADS_n <= #1 1'b0; $display(";A 2930");		//(= P1_P2_P3_ADS_n    0b0)) ;2930
                        P1_P2_P3_State <= #1 3'sb011; $display(";A 2931");		//(= P1_P2_P3_State    0b011)) ;2931
                    end
                3'b011 :
                    begin
                        $display(";A 2932");		//(= P1_P2_P3_State    0b011)) ;2932
                        if ((((P1_P2_P3_READY_n == 1'b0) & (P1_P2_P3_HOLD == 1'b0)) & (P1_P2_P3_RequestPending == 1'b1))) begin
                            $display(";A 2933");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b1))   0b1)) ;2933
                            P1_P2_P3_State <= #1 3'sb010; $display(";A 2935");		//(= P1_P2_P3_State    0b010)) ;2935
                        end
                        else begin
                            $display(";A 2934");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b1))   0b0)) ;2934
                            if (((P1_P2_P3_READY_n == 1'b1) & (P1_P2_P3_NA_n == 1'b1))) begin
                                $display(";A 2936");		//(= (bv-and (bv-comp P1_P2_P3_READY_n  0b1) (bv-comp P1_P2_P3_NA_n  0b1))   0b1)) ;2936
                            end
                            else begin
                                $display(";A 2937");		//(= (bv-and (bv-comp P1_P2_P3_READY_n  0b1) (bv-comp P1_P2_P3_NA_n  0b1))   0b0)) ;2937
                                if ((((P1_P2_P3_RequestPending == 1'b1) | (P1_P2_P3_HOLD == 1'b1)) & ((P1_P2_P3_READY_n == 1'b1) & (P1_P2_P3_NA_n == 1'b0)))) begin
                                    $display(";A 2938");		//(= (bv-and (bv-or (bv-comp P1_P2_P3_RequestPending  0b1) (bv-comp P1_P2_P3_HOLD  0b1)) (bv-and (bv-comp P1_P2_P3_READY_n  0b1) (bv-comp P1_P2_P3_NA_n  0b0)))   0b1)) ;2938
                                    P1_P2_P3_State <= #1 3'sb111; $display(";A 2940");		//(= P1_P2_P3_State    0b111)) ;2940
                                end
                                else begin
                                    $display(";A 2939");		//(= (bv-and (bv-or (bv-comp P1_P2_P3_RequestPending  0b1) (bv-comp P1_P2_P3_HOLD  0b1)) (bv-and (bv-comp P1_P2_P3_READY_n  0b1) (bv-comp P1_P2_P3_NA_n  0b0)))   0b0)) ;2939
                                    if (((((P1_P2_P3_RequestPending == 1'b1) & (P1_P2_P3_HOLD == 1'b0)) & (P1_P2_P3_READY_n == 1'b1)) & (P1_P2_P3_NA_n == 1'b0))) begin
                                        $display(";A 2941");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P2_P3_RequestPending  0b1) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_READY_n  0b1)) (bv-comp P1_P2_P3_NA_n  0b0))   0b1)) ;2941
                                        P1_P2_P3_State <= #1 3'sb110; $display(";A 2943");		//(= P1_P2_P3_State    0b110)) ;2943
                                    end
                                    else begin
                                        $display(";A 2942");		//(= (bv-and (bv-and (bv-and (bv-comp P1_P2_P3_RequestPending  0b1) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_READY_n  0b1)) (bv-comp P1_P2_P3_NA_n  0b0))   0b0)) ;2942
                                        if ((((P1_P2_P3_RequestPending == 1'b0) & (P1_P2_P3_HOLD == 1'b0)) & (P1_P2_P3_READY_n == 1'b0))) begin
                                            $display(";A 2944");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_RequestPending  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_READY_n  0b0))   0b1)) ;2944
                                            P1_P2_P3_State <= #1 3'sb001; $display(";A 2946");		//(= P1_P2_P3_State    0b001)) ;2946
                                        end
                                        else begin
                                            $display(";A 2945");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_RequestPending  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_READY_n  0b0))   0b0)) ;2945
                                            if (((P1_P2_P3_HOLD == 1'b1) & (P1_P2_P3_READY_n == 1'b1))) begin
                                                $display(";A 2947");		//(= (bv-and (bv-comp P1_P2_P3_HOLD  0b1) (bv-comp P1_P2_P3_READY_n  0b1))   0b1)) ;2947
                                                P1_P2_P3_State <= #1 3'sb101; $display(";A 2949");		//(= P1_P2_P3_State    0b101)) ;2949
                                            end
                                            else begin
                                                $display(";A 2948");		//(= (bv-and (bv-comp P1_P2_P3_HOLD  0b1) (bv-comp P1_P2_P3_READY_n  0b1))   0b0)) ;2948
                                                P1_P2_P3_State <= #1 3'sb011; $display(";A 2950");		//(= P1_P2_P3_State    0b011)) ;2950
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P1_P2_P3_StateBS16 <= #1 P1_P2_P3_BS16_n; $display(";A 2951");		//(= P1_P2_P3_StateBS16    P1_P2_P3_BS16_n )) ;2951
                        if ((P1_P2_P3_BS16_n == 1'b0)) begin
                            $display(";A 2952");		//(= (bv-comp P1_P2_P3_BS16_n  0b0)   0b1)) ;2952
                            P1_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 2954");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000001)) ;2954
                        end
                        else begin
                            $display(";A 2953");		//(= (bv-comp P1_P2_P3_BS16_n  0b0)   0b0)) ;2953
                            P1_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 2955");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;2955
                        end
                        P1_P2_P3_StateNA <= #1 P1_P2_P3_NA_n; $display(";A 2956");		//(= P1_P2_P3_StateNA    P1_P2_P3_NA_n )) ;2956
                        P1_P2_P3_ADS_n <= #1 1'b1; $display(";A 2957");		//(= P1_P2_P3_ADS_n    0b1)) ;2957
                    end
                3'b100 :
                    begin
                        $display(";A 2958");		//(= P1_P2_P3_State    0b100)) ;2958
                        if ((((P1_P2_P3_NA_n == 1'b0) & (P1_P2_P3_HOLD == 1'b0)) & (P1_P2_P3_RequestPending == 1'b1))) begin
                            $display(";A 2959");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_NA_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b1))   0b1)) ;2959
                            P1_P2_P3_State <= #1 3'sb110; $display(";A 2961");		//(= P1_P2_P3_State    0b110)) ;2961
                        end
                        else begin
                            $display(";A 2960");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_NA_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b1))   0b0)) ;2960
                            if (((P1_P2_P3_NA_n == 1'b0) & ((P1_P2_P3_HOLD == 1'b1) | (P1_P2_P3_RequestPending == 1'b0)))) begin
                                $display(";A 2962");		//(= (bv-and (bv-comp P1_P2_P3_NA_n  0b0) (bv-or (bv-comp P1_P2_P3_HOLD  0b1) (bv-comp P1_P2_P3_RequestPending  0b0)))   0b1)) ;2962
                                P1_P2_P3_State <= #1 3'sb111; $display(";A 2964");		//(= P1_P2_P3_State    0b111)) ;2964
                            end
                            else begin
                                $display(";A 2963");		//(= (bv-and (bv-comp P1_P2_P3_NA_n  0b0) (bv-or (bv-comp P1_P2_P3_HOLD  0b1) (bv-comp P1_P2_P3_RequestPending  0b0)))   0b0)) ;2963
                                if ((P1_P2_P3_NA_n == 1'b1)) begin
                                    $display(";A 2965");		//(= (bv-comp P1_P2_P3_NA_n  0b1)   0b1)) ;2965
                                    P1_P2_P3_State <= #1 3'sb011; $display(";A 2967");		//(= P1_P2_P3_State    0b011)) ;2967
                                end
                                else begin
                                    $display(";A 2966");		//(= (bv-comp P1_P2_P3_NA_n  0b1)   0b0)) ;2966
                                    P1_P2_P3_State <= #1 3'sb100; $display(";A 2968");		//(= P1_P2_P3_State    0b100)) ;2968
                                end
                            end
                        end
                        P1_P2_P3_StateBS16 <= #1 P1_P2_P3_BS16_n; $display(";A 2969");		//(= P1_P2_P3_StateBS16    P1_P2_P3_BS16_n )) ;2969
                        if ((P1_P2_P3_BS16_n == 1'b0)) begin
                            $display(";A 2970");		//(= (bv-comp P1_P2_P3_BS16_n  0b0)   0b1)) ;2970
                            P1_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 2972");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000001)) ;2972
                        end
                        else begin
                            $display(";A 2971");		//(= (bv-comp P1_P2_P3_BS16_n  0b0)   0b0)) ;2971
                            P1_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 2973");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;2973
                        end
                        P1_P2_P3_StateNA <= #1 P1_P2_P3_NA_n; $display(";A 2974");		//(= P1_P2_P3_StateNA    P1_P2_P3_NA_n )) ;2974
                        P1_P2_P3_ADS_n <= #1 1'b1; $display(";A 2975");		//(= P1_P2_P3_ADS_n    0b1)) ;2975
                    end
                3'b101 :
                    begin
                        $display(";A 2976");		//(= P1_P2_P3_State    0b101)) ;2976
                        if (((P1_P2_P3_HOLD == 1'b0) & (P1_P2_P3_RequestPending == 1'b1))) begin
                            $display(";A 2977");		//(= (bv-and (bv-comp P1_P2_P3_HOLD  0b0) (bv-comp P1_P2_P3_RequestPending  0b1))   0b1)) ;2977
                            P1_P2_P3_State <= #1 3'sb010; $display(";A 2979");		//(= P1_P2_P3_State    0b010)) ;2979
                        end
                        else begin
                            $display(";A 2978");		//(= (bv-and (bv-comp P1_P2_P3_HOLD  0b0) (bv-comp P1_P2_P3_RequestPending  0b1))   0b0)) ;2978
                            if (((P1_P2_P3_HOLD == 1'b0) & (P1_P2_P3_RequestPending == 1'b0))) begin
                                $display(";A 2980");		//(= (bv-and (bv-comp P1_P2_P3_HOLD  0b0) (bv-comp P1_P2_P3_RequestPending  0b0))   0b1)) ;2980
                                P1_P2_P3_State <= #1 3'sb001; $display(";A 2982");		//(= P1_P2_P3_State    0b001)) ;2982
                            end
                            else begin
                                $display(";A 2981");		//(= (bv-and (bv-comp P1_P2_P3_HOLD  0b0) (bv-comp P1_P2_P3_RequestPending  0b0))   0b0)) ;2981
                                P1_P2_P3_State <= #1 3'sb101; $display(";A 2983");		//(= P1_P2_P3_State    0b101)) ;2983
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 2984");		//(= P1_P2_P3_State    0b110)) ;2984
                        P1_P2_P3_Address <= #1 ((P1_P2_P3_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 2985");		//(= P1_P2_P3_Address    (bv-smod (bv-sdiv P1_P2_P3_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;2985
                        P1_P2_P3_BE_n <= #1 P1_P2_P3_ByteEnable; $display(";A 2986");		//(= P1_P2_P3_BE_n    P1_P2_P3_ByteEnable )) ;2986
                        P1_P2_P3_M_IO_n <= #1 P1_P2_P3_MemoryFetch; $display(";A 2987");		//(= P1_P2_P3_M_IO_n    P1_P2_P3_MemoryFetch )) ;2987
                        if ((P1_P2_P3_ReadRequest == 1'b1)) begin
                            $display(";A 2988");		//(= (bv-comp P1_P2_P3_ReadRequest  0b1)   0b1)) ;2988
                            P1_P2_P3_W_R_n <= #1 1'b0; $display(";A 2990");		//(= P1_P2_P3_W_R_n    0b0)) ;2990
                        end
                        else begin
                            $display(";A 2989");		//(= (bv-comp P1_P2_P3_ReadRequest  0b1)   0b0)) ;2989
                            P1_P2_P3_W_R_n <= #1 1'b1; $display(";A 2991");		//(= P1_P2_P3_W_R_n    0b1)) ;2991
                        end
                        if ((P1_P2_P3_CodeFetch == 1'b1)) begin
                            $display(";A 2992");		//(= (bv-comp P1_P2_P3_CodeFetch  0b1)   0b1)) ;2992
                            P1_P2_P3_D_C_n <= #1 1'b0; $display(";A 2994");		//(= P1_P2_P3_D_C_n    0b0)) ;2994
                        end
                        else begin
                            $display(";A 2993");		//(= (bv-comp P1_P2_P3_CodeFetch  0b1)   0b0)) ;2993
                            P1_P2_P3_D_C_n <= #1 1'b1; $display(";A 2995");		//(= P1_P2_P3_D_C_n    0b1)) ;2995
                        end
                        P1_P2_P3_ADS_n <= #1 1'b0; $display(";A 2996");		//(= P1_P2_P3_ADS_n    0b0)) ;2996
                        if ((P1_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 2997");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;2997
                            P1_P2_P3_State <= #1 3'sb100; $display(";A 2999");		//(= P1_P2_P3_State    0b100)) ;2999
                        end
                        else begin
                            $display(";A 2998");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;2998
                            P1_P2_P3_State <= #1 3'sb110; $display(";A 3000");		//(= P1_P2_P3_State    0b110)) ;3000
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 3001");		//(= P1_P2_P3_State    0b111)) ;3001
                        if ((((P1_P2_P3_READY_n == 1'b1) & (P1_P2_P3_RequestPending == 1'b1)) & (P1_P2_P3_HOLD == 1'b0))) begin
                            $display(";A 3002");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b1) (bv-comp P1_P2_P3_RequestPending  0b1)) (bv-comp P1_P2_P3_HOLD  0b0))   0b1)) ;3002
                            P1_P2_P3_State <= #1 3'sb110; $display(";A 3004");		//(= P1_P2_P3_State    0b110)) ;3004
                        end
                        else begin
                            $display(";A 3003");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b1) (bv-comp P1_P2_P3_RequestPending  0b1)) (bv-comp P1_P2_P3_HOLD  0b0))   0b0)) ;3003
                            if (((P1_P2_P3_READY_n == 1'b0) & (P1_P2_P3_HOLD == 1'b1))) begin
                                $display(";A 3005");		//(= (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b1))   0b1)) ;3005
                                P1_P2_P3_State <= #1 3'sb101; $display(";A 3007");		//(= P1_P2_P3_State    0b101)) ;3007
                            end
                            else begin
                                $display(";A 3006");		//(= (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b1))   0b0)) ;3006
                                if ((((P1_P2_P3_READY_n == 1'b0) & (P1_P2_P3_HOLD == 1'b0)) & (P1_P2_P3_RequestPending == 1'b1))) begin
                                    $display(";A 3008");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b1))   0b1)) ;3008
                                    P1_P2_P3_State <= #1 3'sb010; $display(";A 3010");		//(= P1_P2_P3_State    0b010)) ;3010
                                end
                                else begin
                                    $display(";A 3009");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b1))   0b0)) ;3009
                                    if ((((P1_P2_P3_READY_n == 1'b0) & (P1_P2_P3_HOLD == 1'b0)) & (P1_P2_P3_RequestPending == 1'b0))) begin
                                        $display(";A 3011");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b0))   0b1)) ;3011
                                        P1_P2_P3_State <= #1 3'sb001; $display(";A 3013");		//(= P1_P2_P3_State    0b001)) ;3013
                                    end
                                    else begin
                                        $display(";A 3012");		//(= (bv-and (bv-and (bv-comp P1_P2_P3_READY_n  0b0) (bv-comp P1_P2_P3_HOLD  0b0)) (bv-comp P1_P2_P3_RequestPending  0b0))   0b0)) ;3012
                                        P1_P2_P3_State <= #1 3'sb111; $display(";A 3014");		//(= P1_P2_P3_State    0b111)) ;3014
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:4501
    always @(posedge P1_P2_P3_RESET or posedge P1_P2_P3_CLOCK) begin
        if ((P1_P2_P3_RESET == 1'b1)) begin
            $display(";A 3015");		//(= (bv-comp P1_P2_P3_RESET  0b1)   0b1)) ;3015
            P1_P2_P3_State2 = 4'sb0000; $display(";A 3017");		//(= P1_P2_P3_State2    0b0000)) ;3017
            P1_P2_P3_InstQueue[0] = 8'b00000000; $display(";A 3018");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3018
            P1_P2_P3_InstQueue[1] = 8'b00000000; $display(";A 3019");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3019
            P1_P2_P3_InstQueue[2] = 8'b00000000; $display(";A 3020");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3020
            P1_P2_P3_InstQueue[3] = 8'b00000000; $display(";A 3021");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3021
            P1_P2_P3_InstQueue[4] = 8'b00000000; $display(";A 3022");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3022
            P1_P2_P3_InstQueue[5] = 8'b00000000; $display(";A 3023");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3023
            P1_P2_P3_InstQueue[6] = 8'b00000000; $display(";A 3024");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3024
            P1_P2_P3_InstQueue[7] = 8'b00000000; $display(";A 3025");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3025
            P1_P2_P3_InstQueue[8] = 8'b00000000; $display(";A 3026");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3026
            P1_P2_P3_InstQueue[9] = 8'b00000000; $display(";A 3027");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3027
            P1_P2_P3_InstQueue[10] = 8'b00000000; $display(";A 3028");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3028
            P1_P2_P3_InstQueue[11] = 8'b00000000; $display(";A 3029");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3029
            P1_P2_P3_InstQueue[12] = 8'b00000000; $display(";A 3030");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3030
            P1_P2_P3_InstQueue[13] = 8'b00000000; $display(";A 3031");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3031
            P1_P2_P3_InstQueue[14] = 8'b00000000; $display(";A 3032");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3032
            P1_P2_P3_InstQueue[15] = 8'b00000000; $display(";A 3033");		//(= P1_P2_P3_InstQueue    0b00000000)) ;3033
            P1_P2_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 3034");		//(= P1_P2_P3_InstQueueRd_Addr    0b00000)) ;3034
            P1_P2_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 3035");		//(= P1_P2_P3_InstQueueWr_Addr    0b00000)) ;3035
            P1_P2_P3_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 3036");		//(= P1_P2_P3_InstAddrPointer    0b00000000000000000000000000000000)) ;3036
            P1_P2_P3_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 3037");		//(= P1_P2_P3_PhyAddrPointer    0b00000000000000000000000000000000)) ;3037
            P1_P2_P3_Extended = 1'b0; $display(";A 3038");		//(= P1_P2_P3_Extended    0b0)) ;3038
            P1_P2_P3_More = 1'b0; $display(";A 3039");		//(= P1_P2_P3_More    0b0)) ;3039
            P1_P2_P3_Flush = 1'b0; $display(";A 3040");		//(= P1_P2_P3_Flush    0b0)) ;3040
            P1_P2_P3_lWord = 16'sb0000000000000000; $display(";A 3041");		//(= P1_P2_P3_lWord    0b0000000000000000)) ;3041
            P1_P2_P3_uWord = 15'sb000000000000000; $display(";A 3042");		//(= P1_P2_P3_uWord    0b000000000000000)) ;3042
            P1_P2_P3_fWord = 32'sb00000000000000000000000000000000; $display(";A 3043");		//(= P1_P2_P3_fWord    0b00000000000000000000000000000000)) ;3043
            P1_P2_P3_CodeFetch <= #1 1'b0; $display(";A 3044");		//(= P1_P2_P3_CodeFetch    0b0)) ;3044
            P1_P2_P3_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 3045");		//(= P1_P2_P3_Datao    0b00000000000000000000000000000000)) ;3045
            P1_P2_P3_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 3046");		//(= P1_P2_P3_EAX    0b00000000000000000000000000000000)) ;3046
            P1_P2_P3_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 3047");		//(= P1_P2_P3_EBX    0b00000000000000000000000000000000)) ;3047
            P1_P2_P3_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 3048");		//(= P1_P2_P3_rEIP    0b00000000000000000000000000000000)) ;3048
            P1_P2_P3_ReadRequest <= #1 1'b0; $display(";A 3049");		//(= P1_P2_P3_ReadRequest    0b0)) ;3049
            P1_P2_P3_MemoryFetch <= #1 1'b0; $display(";A 3050");		//(= P1_P2_P3_MemoryFetch    0b0)) ;3050
            P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3051");		//(= P1_P2_P3_RequestPending    0b0)) ;3051
        end
        else begin
            $display(";A 3016");		//(= (bv-comp P1_P2_P3_RESET  0b1)   0b0)) ;3016
            case (P1_P2_P3_State2)
                4'b0000 :
                    begin
                        $display(";A 3052");		//(= P1_P2_P3_State2    0b0000)) ;3052
                        P1_P2_P3_PhyAddrPointer = P1_P2_P3_rEIP; $display(";A 3053");		//(= P1_P2_P3_PhyAddrPointer    P1_P2_P3_rEIP )) ;3053
                        P1_P2_P3_InstAddrPointer = P1_P2_P3_PhyAddrPointer; $display(";A 3054");		//(= P1_P2_P3_InstAddrPointer    P1_P2_P3_PhyAddrPointer )) ;3054
                        P1_P2_P3_State2 = 4'sb0001; $display(";A 3055");		//(= P1_P2_P3_State2    0b0001)) ;3055
                        P1_P2_P3_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 3056");		//(= P1_P2_P3_rEIP    0b00000000000011111111111111110000)) ;3056
                        P1_P2_P3_ReadRequest <= #1 1'b1; $display(";A 3057");		//(= P1_P2_P3_ReadRequest    0b1)) ;3057
                        P1_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 3058");		//(= P1_P2_P3_MemoryFetch    0b1)) ;3058
                        P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3059");		//(= P1_P2_P3_RequestPending    0b1)) ;3059
                    end
                4'b0001 :
                    begin
                        $display(";A 3060");		//(= P1_P2_P3_State2    0b0001)) ;3060
                        P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3061");		//(= P1_P2_P3_RequestPending    0b1)) ;3061
                        P1_P2_P3_ReadRequest <= #1 1'b1; $display(";A 3062");		//(= P1_P2_P3_ReadRequest    0b1)) ;3062
                        P1_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 3063");		//(= P1_P2_P3_MemoryFetch    0b1)) ;3063
                        P1_P2_P3_CodeFetch <= #1 1'b1; $display(";A 3064");		//(= P1_P2_P3_CodeFetch    0b1)) ;3064
                        if ((P1_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 3065");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3065
                            P1_P2_P3_State2 = 4'sb0010; $display(";A 3067");		//(= P1_P2_P3_State2    0b0010)) ;3067
                        end
                        else begin
                            $display(";A 3066");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3066
                            P1_P2_P3_State2 = 4'sb0001; $display(";A 3068");		//(= P1_P2_P3_State2    0b0001)) ;3068
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 3069");		//(= P1_P2_P3_State2    0b0010)) ;3069
                        P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3070");		//(= P1_P2_P3_RequestPending    0b0)) ;3070
                        P1_P2_P3_InstQueue[P1_P2_P3_InstQueueWr_Addr] = (P1_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 3071");		//(= P1_P2_P3_InstQueue    (bv-smod P1_P2_P3_Datai  0b00000000000000000000000100000000))) ;3071
                        P1_P2_P3_InstQueueWr_Addr = ((P1_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3072");		//(= P1_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3072
                        P1_P2_P3_InstQueue[P1_P2_P3_InstQueueWr_Addr] = (P1_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 3073");		//(= P1_P2_P3_InstQueue    (bv-smod P1_P2_P3_Datai  0b00000000000000000000000100000000))) ;3073
                        P1_P2_P3_InstQueueWr_Addr = ((P1_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3074");		//(= P1_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3074
                        if ((P1_P2_P3_StateBS16 == 1'b1)) begin
                            $display(";A 3075");		//(= (bv-comp P1_P2_P3_StateBS16  0b1)   0b1)) ;3075
                            P1_P2_P3_InstQueue[P1_P2_P3_InstQueueWr_Addr] = ((P1_P2_P3_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 3077");		//(= P1_P2_P3_InstQueue    (bv-smod (bv-sdiv P1_P2_P3_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;3077
                            P1_P2_P3_InstQueueWr_Addr = ((P1_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3078");		//(= P1_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3078
                            P1_P2_P3_InstQueue[P1_P2_P3_InstQueueWr_Addr] = ((P1_P2_P3_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 3079");		//(= P1_P2_P3_InstQueue    (bv-smod (bv-sdiv P1_P2_P3_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;3079
                            P1_P2_P3_InstQueueWr_Addr = ((P1_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3080");		//(= P1_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3080
                            P1_P2_P3_PhyAddrPointer = (P1_P2_P3_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 3081");		//(= P1_P2_P3_PhyAddrPointer    (bv-add P1_P2_P3_PhyAddrPointer  0b00000000000000000000000000000100))) ;3081
                            P1_P2_P3_State2 = 4'sb0101; $display(";A 3082");		//(= P1_P2_P3_State2    0b0101)) ;3082
                        end
                        else begin
                            $display(";A 3076");		//(= (bv-comp P1_P2_P3_StateBS16  0b1)   0b0)) ;3076
                            P1_P2_P3_PhyAddrPointer = (P1_P2_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3083");		//(= P1_P2_P3_PhyAddrPointer    (bv-add P1_P2_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;3083
                            if ((P1_P2_P3_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 3084");		//(= (bool-to-bv (bv-slt P1_P2_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;3084
                                P1_P2_P3_rEIP <= #1 (-P1_P2_P3_PhyAddrPointer); $display(";A 3086");		//(= P1_P2_P3_rEIP    (bv-neg P1_P2_P3_PhyAddrPointer ))) ;3086
                            end
                            else begin
                                $display(";A 3085");		//(= (bool-to-bv (bv-slt P1_P2_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;3085
                                P1_P2_P3_rEIP <= #1 P1_P2_P3_PhyAddrPointer; $display(";A 3087");		//(= P1_P2_P3_rEIP    P1_P2_P3_PhyAddrPointer )) ;3087
                            end
                            P1_P2_P3_State2 = 4'sb0011; $display(";A 3088");		//(= P1_P2_P3_State2    0b0011)) ;3088
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 3089");		//(= P1_P2_P3_State2    0b0011)) ;3089
                        P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3090");		//(= P1_P2_P3_RequestPending    0b1)) ;3090
                        if ((P1_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 3091");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3091
                            P1_P2_P3_State2 = 4'sb0100; $display(";A 3093");		//(= P1_P2_P3_State2    0b0100)) ;3093
                        end
                        else begin
                            $display(";A 3092");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3092
                            P1_P2_P3_State2 = 4'sb0011; $display(";A 3094");		//(= P1_P2_P3_State2    0b0011)) ;3094
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 3095");		//(= P1_P2_P3_State2    0b0100)) ;3095
                        P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3096");		//(= P1_P2_P3_RequestPending    0b0)) ;3096
                        P1_P2_P3_InstQueue[P1_P2_P3_InstQueueWr_Addr] = (P1_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 3097");		//(= P1_P2_P3_InstQueue    (bv-smod P1_P2_P3_Datai  0b00000000000000000000000100000000))) ;3097
                        P1_P2_P3_InstQueueWr_Addr = ((P1_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3098");		//(= P1_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3098
                        P1_P2_P3_InstQueue[P1_P2_P3_InstQueueWr_Addr] = (P1_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 3099");		//(= P1_P2_P3_InstQueue    (bv-smod P1_P2_P3_Datai  0b00000000000000000000000100000000))) ;3099
                        P1_P2_P3_InstQueueWr_Addr = ((P1_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3100");		//(= P1_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3100
                        P1_P2_P3_PhyAddrPointer = (P1_P2_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3101");		//(= P1_P2_P3_PhyAddrPointer    (bv-add P1_P2_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;3101
                        P1_P2_P3_State2 = 4'sb0101; $display(";A 3102");		//(= P1_P2_P3_State2    0b0101)) ;3102
                    end
                4'b0101 :
                    begin
                        $display(";A 3103");		//(= P1_P2_P3_State2    0b0101)) ;3103
                        case (P1_P2_P3_InstQueue[P1_P2_P3_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 3104");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b10010000)) ;3104
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3105");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3105
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3106");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3106
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3107");		//(= P1_P2_P3_Flush    0b0)) ;3107
                                    P1_P2_P3_More = 1'b0; $display(";A 3108");		//(= P1_P2_P3_More    0b0)) ;3108
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 3109");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b01100110)) ;3109
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3110");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3110
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3111");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3111
                                    P1_P2_P3_Extended = 1'b1; $display(";A 3112");		//(= P1_P2_P3_Extended    0b1)) ;3112
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3113");		//(= P1_P2_P3_Flush    0b0)) ;3113
                                    P1_P2_P3_More = 1'b0; $display(";A 3114");		//(= P1_P2_P3_More    0b0)) ;3114
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 3115");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b11101011)) ;3115
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 3116");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;3116
                                        if ((P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 3118");		//(= (bool-to-bv (bv-gt P1_P2_P3_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;3118
                                            P1_P2_P3_PhyAddrPointer = ((P1_P2_P3_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 3120");		//(= P1_P2_P3_PhyAddrPointer    (bv-sub (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P1_P2_P3_InstQueue 0 )))) ;3120
                                            P1_P2_P3_InstAddrPointer = P1_P2_P3_PhyAddrPointer; $display(";A 3121");		//(= P1_P2_P3_InstAddrPointer    P1_P2_P3_PhyAddrPointer )) ;3121
                                        end
                                        else begin
                                            $display(";A 3119");		//(= (bool-to-bv (bv-gt P1_P2_P3_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;3119
                                            P1_P2_P3_PhyAddrPointer = ((P1_P2_P3_InstAddrPointer + 32'b00000000000000000000000000000010) + P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 3122");		//(= P1_P2_P3_PhyAddrPointer    (bv-add (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000010) P1_P2_P3_InstQueue 0 ))) ;3122
                                            P1_P2_P3_InstAddrPointer = P1_P2_P3_PhyAddrPointer; $display(";A 3123");		//(= P1_P2_P3_InstAddrPointer    P1_P2_P3_PhyAddrPointer )) ;3123
                                        end
                                        P1_P2_P3_Flush = 1'b1; $display(";A 3124");		//(= P1_P2_P3_Flush    0b1)) ;3124
                                        P1_P2_P3_More = 1'b0; $display(";A 3125");		//(= P1_P2_P3_More    0b0)) ;3125
                                    end
                                    else begin
                                        $display(";A 3117");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;3117
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3126");		//(= P1_P2_P3_Flush    0b0)) ;3126
                                        P1_P2_P3_More = 1'b1; $display(";A 3127");		//(= P1_P2_P3_More    0b1)) ;3127
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 3128");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b11101001)) ;3128
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 3129");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;3129
                                        P1_P2_P3_PhyAddrPointer = ((P1_P2_P3_InstAddrPointer + 32'b00000000000000000000000000000101) + P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 3131");		//(= P1_P2_P3_PhyAddrPointer    (bv-add (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000101) P1_P2_P3_InstQueue 0 ))) ;3131
                                        P1_P2_P3_InstAddrPointer = P1_P2_P3_PhyAddrPointer; $display(";A 3132");		//(= P1_P2_P3_InstAddrPointer    P1_P2_P3_PhyAddrPointer )) ;3132
                                        P1_P2_P3_Flush = 1'b1; $display(";A 3133");		//(= P1_P2_P3_Flush    0b1)) ;3133
                                        P1_P2_P3_More = 1'b0; $display(";A 3134");		//(= P1_P2_P3_More    0b0)) ;3134
                                    end
                                    else begin
                                        $display(";A 3130");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;3130
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3135");		//(= P1_P2_P3_Flush    0b0)) ;3135
                                        P1_P2_P3_More = 1'b1; $display(";A 3136");		//(= P1_P2_P3_More    0b1)) ;3136
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 3137");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b11101010)) ;3137
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3138");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3138
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3139");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3139
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3140");		//(= P1_P2_P3_Flush    0b0)) ;3140
                                    P1_P2_P3_More = 1'b0; $display(";A 3141");		//(= P1_P2_P3_More    0b0)) ;3141
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 3142");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b10110000)) ;3142
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3143");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3143
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3144");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3144
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3145");		//(= P1_P2_P3_Flush    0b0)) ;3145
                                    P1_P2_P3_More = 1'b0; $display(";A 3146");		//(= P1_P2_P3_More    0b0)) ;3146
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 3147");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b10111000)) ;3147
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 3148");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;3148
                                        P1_P2_P3_EAX <= #1 ((((P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 3150");		//(= P1_P2_P3_EAX    (bv-add (bv-add (bv-add (bv-mul P1_P2_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P2_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P2_P3_InstQueue 0  0b00000000000000000000000100000000)) P1_P2_P3_InstQueue 0 ))) ;3150
                                        P1_P2_P3_More = 1'b0; $display(";A 3151");		//(= P1_P2_P3_More    0b0)) ;3151
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3152");		//(= P1_P2_P3_Flush    0b0)) ;3152
                                        P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 3153");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;3153
                                        P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 3154");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;3154
                                    end
                                    else begin
                                        $display(";A 3149");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;3149
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3155");		//(= P1_P2_P3_Flush    0b0)) ;3155
                                        P1_P2_P3_More = 1'b1; $display(";A 3156");		//(= P1_P2_P3_More    0b1)) ;3156
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 3157");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b10111011)) ;3157
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 3158");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;3158
                                        P1_P2_P3_EBX <= #1 ((((P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P1_P2_P3_InstQueue[((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 3160");		//(= P1_P2_P3_EBX    (bv-add (bv-add (bv-add (bv-mul P1_P2_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P1_P2_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P1_P2_P3_InstQueue 0  0b00000000000000000000000100000000)) P1_P2_P3_InstQueue 0 ))) ;3160
                                        P1_P2_P3_More = 1'b0; $display(";A 3161");		//(= P1_P2_P3_More    0b0)) ;3161
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3162");		//(= P1_P2_P3_Flush    0b0)) ;3162
                                        P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 3163");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;3163
                                        P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 3164");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;3164
                                    end
                                    else begin
                                        $display(";A 3159");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;3159
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3165");		//(= P1_P2_P3_Flush    0b0)) ;3165
                                        P1_P2_P3_More = 1'b1; $display(";A 3166");		//(= P1_P2_P3_More    0b1)) ;3166
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 3167");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b10001011)) ;3167
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 3168");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;3168
                                        if ((P1_P2_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 3170");		//(= (bool-to-bv (bv-slt P1_P2_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;3170
                                            P1_P2_P3_rEIP <= #1 (-P1_P2_P3_EBX); $display(";A 3172");		//(= P1_P2_P3_rEIP    (bv-neg P1_P2_P3_EBX ))) ;3172
                                        end
                                        else begin
                                            $display(";A 3171");		//(= (bool-to-bv (bv-slt P1_P2_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;3171
                                            P1_P2_P3_rEIP <= #1 P1_P2_P3_EBX; $display(";A 3173");		//(= P1_P2_P3_rEIP    P1_P2_P3_EBX )) ;3173
                                        end
                                        P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3174");		//(= P1_P2_P3_RequestPending    0b1)) ;3174
                                        P1_P2_P3_ReadRequest <= #1 1'b1; $display(";A 3175");		//(= P1_P2_P3_ReadRequest    0b1)) ;3175
                                        P1_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 3176");		//(= P1_P2_P3_MemoryFetch    0b1)) ;3176
                                        P1_P2_P3_CodeFetch <= #1 1'b0; $display(";A 3177");		//(= P1_P2_P3_CodeFetch    0b0)) ;3177
                                        if ((P1_P2_P3_READY_n == 1'b0)) begin
                                            $display(";A 3178");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3178
                                            P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3180");		//(= P1_P2_P3_RequestPending    0b0)) ;3180
                                            P1_P2_P3_uWord = (P1_P2_P3_Datai % 32'b00000000000000001000000000000000); $display(";A 3181");		//(= P1_P2_P3_uWord    (bv-smod P1_P2_P3_Datai  0b00000000000000001000000000000000))) ;3181
                                            if ((P1_P2_P3_StateBS16 == 1'b1)) begin
                                                $display(";A 3182");		//(= (bv-comp P1_P2_P3_StateBS16  0b1)   0b1)) ;3182
                                                P1_P2_P3_lWord = (P1_P2_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 3184");		//(= P1_P2_P3_lWord    (bv-smod P1_P2_P3_Datai  0b00000000000000010000000000000000))) ;3184
                                            end
                                            else begin
                                                $display(";A 3183");		//(= (bv-comp P1_P2_P3_StateBS16  0b1)   0b0)) ;3183
                                                P1_P2_P3_rEIP <= #1 (P1_P2_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 3185");		//(= P1_P2_P3_rEIP    (bv-add P1_P2_P3_rEIP  0b00000000000000000000000000000010))) ;3185
                                                P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3186");		//(= P1_P2_P3_RequestPending    0b1)) ;3186
                                                if ((P1_P2_P3_READY_n == 1'b0)) begin
                                                    $display(";A 3187");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3187
                                                    P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3189");		//(= P1_P2_P3_RequestPending    0b0)) ;3189
                                                    P1_P2_P3_lWord = (P1_P2_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 3190");		//(= P1_P2_P3_lWord    (bv-smod P1_P2_P3_Datai  0b00000000000000010000000000000000))) ;3190
                                                end
                                                else begin
                                                    $display(";A 3188");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3188
                                                end
                                            end
                                            if ((P1_P2_P3_READY_n == 1'b0)) begin
                                                $display(";A 3191");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3191
                                                P1_P2_P3_EAX <= #1 ((P1_P2_P3_uWord * 32'b00000000000000010000000000000000) + P1_P2_P3_lWord); $display(";A 3193");		//(= P1_P2_P3_EAX    (bv-add (bv-mul P1_P2_P3_uWord  0b00000000000000010000000000000000) P1_P2_P3_lWord ))) ;3193
                                                P1_P2_P3_More = 1'b0; $display(";A 3194");		//(= P1_P2_P3_More    0b0)) ;3194
                                                P1_P2_P3_Flush = 1'b0; $display(";A 3195");		//(= P1_P2_P3_Flush    0b0)) ;3195
                                                P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3196");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;3196
                                                P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 3197");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;3197
                                            end
                                            else begin
                                                $display(";A 3192");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3192
                                            end
                                        end
                                        else begin
                                            $display(";A 3179");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3179
                                        end
                                    end
                                    else begin
                                        $display(";A 3169");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;3169
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3198");		//(= P1_P2_P3_Flush    0b0)) ;3198
                                        P1_P2_P3_More = 1'b1; $display(";A 3199");		//(= P1_P2_P3_More    0b1)) ;3199
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 3200");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b10001001)) ;3200
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 3201");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;3201
                                        if ((P1_P2_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 3203");		//(= (bool-to-bv (bv-slt P1_P2_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;3203
                                            P1_P2_P3_rEIP <= #1 P1_P2_P3_EBX; $display(";A 3205");		//(= P1_P2_P3_rEIP    P1_P2_P3_EBX )) ;3205
                                        end
                                        else begin
                                            $display(";A 3204");		//(= (bool-to-bv (bv-slt P1_P2_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;3204
                                            P1_P2_P3_rEIP <= #1 P1_P2_P3_EBX; $display(";A 3206");		//(= P1_P2_P3_rEIP    P1_P2_P3_EBX )) ;3206
                                        end
                                        P1_P2_P3_lWord = (P1_P2_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 3207");		//(= P1_P2_P3_lWord    (bv-smod P1_P2_P3_EAX  0b00000000000000010000000000000000))) ;3207
                                        P1_P2_P3_uWord = ((P1_P2_P3_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 3208");		//(= P1_P2_P3_uWord    (bv-smod (bv-sdiv P1_P2_P3_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;3208
                                        P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3209");		//(= P1_P2_P3_RequestPending    0b1)) ;3209
                                        P1_P2_P3_ReadRequest <= #1 1'b0; $display(";A 3210");		//(= P1_P2_P3_ReadRequest    0b0)) ;3210
                                        P1_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 3211");		//(= P1_P2_P3_MemoryFetch    0b1)) ;3211
                                        P1_P2_P3_CodeFetch <= #1 1'b0; $display(";A 3212");		//(= P1_P2_P3_CodeFetch    0b0)) ;3212
                                        if (((P1_P2_P3_State == 32'b00000000000000000000000000000010) | (P1_P2_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 3213");		//(= (bv-or (bv-comp P1_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P3_State  0b00000000000000000000000000000100))   0b1)) ;3213
                                            P1_P2_P3_Datao <= #1 ((P1_P2_P3_uWord * 32'b00000000000000010000000000000000) + P1_P2_P3_lWord); $display(";A 3215");		//(= P1_P2_P3_Datao    (bv-add (bv-mul P1_P2_P3_uWord  0b00000000000000010000000000000000) P1_P2_P3_lWord ))) ;3215
                                            if ((P1_P2_P3_READY_n == 1'b0)) begin
                                                $display(";A 3216");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3216
                                                P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3218");		//(= P1_P2_P3_RequestPending    0b0)) ;3218
                                                if ((P1_P2_P3_StateBS16 == 1'b0)) begin
                                                    $display(";A 3219");		//(= (bv-comp P1_P2_P3_StateBS16  0b0)   0b1)) ;3219
                                                    P1_P2_P3_rEIP <= #1 (P1_P2_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 3221");		//(= P1_P2_P3_rEIP    (bv-add P1_P2_P3_rEIP  0b00000000000000000000000000000010))) ;3221
                                                    P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3222");		//(= P1_P2_P3_RequestPending    0b1)) ;3222
                                                    P1_P2_P3_ReadRequest <= #1 1'b0; $display(";A 3223");		//(= P1_P2_P3_ReadRequest    0b0)) ;3223
                                                    P1_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 3224");		//(= P1_P2_P3_MemoryFetch    0b1)) ;3224
                                                    P1_P2_P3_CodeFetch <= #1 1'b0; $display(";A 3225");		//(= P1_P2_P3_CodeFetch    0b0)) ;3225
                                                    P1_P2_P3_State2 = 4'sb0110; $display(";A 3226");		//(= P1_P2_P3_State2    0b0110)) ;3226
                                                end
                                                else begin
                                                    $display(";A 3220");		//(= (bv-comp P1_P2_P3_StateBS16  0b0)   0b0)) ;3220
                                                end
                                                P1_P2_P3_More = 1'b0; $display(";A 3227");		//(= P1_P2_P3_More    0b0)) ;3227
                                                P1_P2_P3_Flush = 1'b0; $display(";A 3228");		//(= P1_P2_P3_Flush    0b0)) ;3228
                                                P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3229");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;3229
                                                P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 3230");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;3230
                                            end
                                            else begin
                                                $display(";A 3217");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3217
                                            end
                                        end
                                        else begin
                                            $display(";A 3214");		//(= (bv-or (bv-comp P1_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P3_State  0b00000000000000000000000000000100))   0b0)) ;3214
                                        end
                                    end
                                    else begin
                                        $display(";A 3202");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;3202
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3231");		//(= P1_P2_P3_Flush    0b0)) ;3231
                                        P1_P2_P3_More = 1'b1; $display(";A 3232");		//(= P1_P2_P3_More    0b1)) ;3232
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 3233");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b11100100)) ;3233
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 3234");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;3234
                                        P1_P2_P3_rEIP <= #1 (P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 3236");		//(= P1_P2_P3_rEIP    (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;3236
                                        P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3237");		//(= P1_P2_P3_RequestPending    0b1)) ;3237
                                        P1_P2_P3_ReadRequest <= #1 1'b1; $display(";A 3238");		//(= P1_P2_P3_ReadRequest    0b1)) ;3238
                                        P1_P2_P3_MemoryFetch <= #1 1'b0; $display(";A 3239");		//(= P1_P2_P3_MemoryFetch    0b0)) ;3239
                                        P1_P2_P3_CodeFetch <= #1 1'b0; $display(";A 3240");		//(= P1_P2_P3_CodeFetch    0b0)) ;3240
                                        if ((P1_P2_P3_READY_n == 1'b0)) begin
                                            $display(";A 3241");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3241
                                            P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3243");		//(= P1_P2_P3_RequestPending    0b0)) ;3243
                                            P1_P2_P3_EAX <= #1 P1_P2_P3_Datai; $display(";A 3244");		//(= P1_P2_P3_EAX    P1_P2_P3_Datai )) ;3244
                                            P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3245");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;3245
                                            P1_P2_P3_InstQueueRd_Addr = (P1_P2_P3_InstQueueRd_Addr + 5'b00010); $display(";A 3246");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-add P1_P2_P3_InstQueueRd_Addr  0b00010))) ;3246
                                            P1_P2_P3_Flush = 1'b0; $display(";A 3247");		//(= P1_P2_P3_Flush    0b0)) ;3247
                                            P1_P2_P3_More = 1'b0; $display(";A 3248");		//(= P1_P2_P3_More    0b0)) ;3248
                                        end
                                        else begin
                                            $display(";A 3242");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3242
                                        end
                                    end
                                    else begin
                                        $display(";A 3235");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;3235
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3249");		//(= P1_P2_P3_Flush    0b0)) ;3249
                                        P1_P2_P3_More = 1'b1; $display(";A 3250");		//(= P1_P2_P3_More    0b1)) ;3250
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 3251");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b11100110)) ;3251
                                    if (((P1_P2_P3_InstQueueWr_Addr - P1_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 3252");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;3252
                                        P1_P2_P3_rEIP <= #1 (P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 3254");		//(= P1_P2_P3_rEIP    (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;3254
                                        P1_P2_P3_RequestPending <= #1 1'b1; $display(";A 3255");		//(= P1_P2_P3_RequestPending    0b1)) ;3255
                                        P1_P2_P3_ReadRequest <= #1 1'b0; $display(";A 3256");		//(= P1_P2_P3_ReadRequest    0b0)) ;3256
                                        P1_P2_P3_MemoryFetch <= #1 1'b0; $display(";A 3257");		//(= P1_P2_P3_MemoryFetch    0b0)) ;3257
                                        P1_P2_P3_CodeFetch <= #1 1'b0; $display(";A 3258");		//(= P1_P2_P3_CodeFetch    0b0)) ;3258
                                        if (((P1_P2_P3_State == 32'b00000000000000000000000000000010) | (P1_P2_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 3259");		//(= (bv-or (bv-comp P1_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P3_State  0b00000000000000000000000000000100))   0b1)) ;3259
                                            P1_P2_P3_fWord = (P1_P2_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 3261");		//(= P1_P2_P3_fWord    (bv-smod P1_P2_P3_EAX  0b00000000000000010000000000000000))) ;3261
                                            P1_P2_P3_Datao <= #1 P1_P2_P3_fWord; $display(";A 3262");		//(= P1_P2_P3_Datao    P1_P2_P3_fWord )) ;3262
                                            if ((P1_P2_P3_READY_n == 1'b0)) begin
                                                $display(";A 3263");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3263
                                                P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3265");		//(= P1_P2_P3_RequestPending    0b0)) ;3265
                                                P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3266");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;3266
                                                P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 3267");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;3267
                                                P1_P2_P3_Flush = 1'b0; $display(";A 3268");		//(= P1_P2_P3_Flush    0b0)) ;3268
                                                P1_P2_P3_More = 1'b0; $display(";A 3269");		//(= P1_P2_P3_More    0b0)) ;3269
                                            end
                                            else begin
                                                $display(";A 3264");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3264
                                            end
                                        end
                                        else begin
                                            $display(";A 3260");		//(= (bv-or (bv-comp P1_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P1_P2_P3_State  0b00000000000000000000000000000100))   0b0)) ;3260
                                        end
                                    end
                                    else begin
                                        $display(";A 3253");		//(= (bool-to-bv (bv-ge (bv-sub P1_P2_P3_InstQueueWr_Addr  P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;3253
                                        P1_P2_P3_Flush = 1'b0; $display(";A 3270");		//(= P1_P2_P3_Flush    0b0)) ;3270
                                        P1_P2_P3_More = 1'b1; $display(";A 3271");		//(= P1_P2_P3_More    0b1)) ;3271
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 3272");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b00000100)) ;3272
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3273");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3273
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3274");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3274
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3275");		//(= P1_P2_P3_Flush    0b0)) ;3275
                                    P1_P2_P3_More = 1'b0; $display(";A 3276");		//(= P1_P2_P3_More    0b0)) ;3276
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 3277");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b00000101)) ;3277
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3278");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3278
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3279");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3279
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3280");		//(= P1_P2_P3_Flush    0b0)) ;3280
                                    P1_P2_P3_More = 1'b0; $display(";A 3281");		//(= P1_P2_P3_More    0b0)) ;3281
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 3282");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b11010000)) ;3282
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3283");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;3283
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 3284");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;3284
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3285");		//(= P1_P2_P3_Flush    0b0)) ;3285
                                    P1_P2_P3_More = 1'b0; $display(";A 3286");		//(= P1_P2_P3_More    0b0)) ;3286
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 3287");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b11000000)) ;3287
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 3288");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;3288
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 3289");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;3289
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3290");		//(= P1_P2_P3_Flush    0b0)) ;3290
                                    P1_P2_P3_More = 1'b0; $display(";A 3291");		//(= P1_P2_P3_More    0b0)) ;3291
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 3292");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b01000000)) ;3292
                                    P1_P2_P3_EAX <= #1 (P1_P2_P3_EAX + 32'sb00000000000000000000000000000001); $display(";A 3293");		//(= P1_P2_P3_EAX    (bv-add P1_P2_P3_EAX  0b00000000000000000000000000000001))) ;3293
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3294");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3294
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3295");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3295
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3296");		//(= P1_P2_P3_Flush    0b0)) ;3296
                                    P1_P2_P3_More = 1'b0; $display(";A 3297");		//(= P1_P2_P3_More    0b0)) ;3297
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 3298");		//(= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr )   0b01000011)) ;3298
                                    P1_P2_P3_EBX <= #1 (P1_P2_P3_EBX + 32'sb00000000000000000000000000000001); $display(";A 3299");		//(= P1_P2_P3_EBX    (bv-add P1_P2_P3_EBX  0b00000000000000000000000000000001))) ;3299
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3300");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3300
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3301");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3301
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3302");		//(= P1_P2_P3_Flush    0b0)) ;3302
                                    P1_P2_P3_More = 1'b0; $display(";A 3303");		//(= P1_P2_P3_More    0b0)) ;3303
                                end
                            default:
                                begin
                                    $display(";A 3304");		//(= (and (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b10010000) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b01100110) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b11101011) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b11101001) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b11101010) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b10110000) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b10111000) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b10111011) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b10001011) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b10001001) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b11100100) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b11100110) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b00000100) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b00000101) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b11010000) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b11000000) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b01000000) (/= ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ) 0b01000011))   true)) ;3304
                                    P1_P2_P3_InstAddrPointer = (P1_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 3305");		//(= P1_P2_P3_InstAddrPointer    (bv-add P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;3305
                                    P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3306");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3306
                                    P1_P2_P3_Flush = 1'b0; $display(";A 3307");		//(= P1_P2_P3_Flush    0b0)) ;3307
                                    P1_P2_P3_More = 1'b0; $display(";A 3308");		//(= P1_P2_P3_More    0b0)) ;3308
                                end
                        endcase
                        if (((~(P1_P2_P3_InstQueueRd_Addr < P1_P2_P3_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P1_P2_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P1_P2_P3_Flush) | P1_P2_P3_More))) begin
                            $display(";A 3309");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P2_P3_InstQueueRd_Addr  P1_P2_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P2_P3_Flush ) P1_P2_P3_More ))   0b1)) ;3309
                            P1_P2_P3_State2 = 4'sb0111; $display(";A 3311");		//(= P1_P2_P3_State2    0b0111)) ;3311
                        end
                        else begin
                            $display(";A 3310");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P1_P2_P3_InstQueueRd_Addr  P1_P2_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P1_P2_P3_Flush ) P1_P2_P3_More ))   0b0)) ;3310
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 3312");		//(= P1_P2_P3_State2    0b0110)) ;3312
                        P1_P2_P3_Datao <= #1 ((P1_P2_P3_uWord * 32'b00000000000000010000000000000000) + P1_P2_P3_lWord); $display(";A 3313");		//(= P1_P2_P3_Datao    (bv-add (bv-mul P1_P2_P3_uWord  0b00000000000000010000000000000000) P1_P2_P3_lWord ))) ;3313
                        if ((P1_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 3314");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b1)) ;3314
                            P1_P2_P3_RequestPending <= #1 1'b0; $display(";A 3316");		//(= P1_P2_P3_RequestPending    0b0)) ;3316
                            P1_P2_P3_State2 = 4'sb0101; $display(";A 3317");		//(= P1_P2_P3_State2    0b0101)) ;3317
                        end
                        else begin
                            $display(";A 3315");		//(= (bv-comp P1_P2_P3_READY_n  0b0)   0b0)) ;3315
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 3318");		//(= P1_P2_P3_State2    0b0111)) ;3318
                        if (P1_P2_P3_Flush) begin
                            $display(";A 3319");		//(= P1_P2_P3_Flush    0b1)) ;3319
                            P1_P2_P3_InstQueueRd_Addr = 5'sb00001; $display(";A 3321");		//(= P1_P2_P3_InstQueueRd_Addr    0b00001)) ;3321
                            P1_P2_P3_InstQueueWr_Addr = 5'sb00001; $display(";A 3322");		//(= P1_P2_P3_InstQueueWr_Addr    0b00001)) ;3322
                            if ((P1_P2_P3_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 3323");		//(= (bool-to-bv (bv-slt P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;3323
                                P1_P2_P3_fWord = (-P1_P2_P3_InstAddrPointer); $display(";A 3325");		//(= P1_P2_P3_fWord    (bv-neg P1_P2_P3_InstAddrPointer ))) ;3325
                            end
                            else begin
                                $display(";A 3324");		//(= (bool-to-bv (bv-slt P1_P2_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;3324
                                P1_P2_P3_fWord = P1_P2_P3_InstAddrPointer; $display(";A 3326");		//(= P1_P2_P3_fWord    P1_P2_P3_InstAddrPointer )) ;3326
                            end
                            if (((P1_P2_P3_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 3327");		//(= (bv-comp (bv-smod P1_P2_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;3327
                                P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + (P1_P2_P3_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 3329");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  (bv-smod P1_P2_P3_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;3329
                            end
                            else begin
                                $display(";A 3328");		//(= (bv-comp (bv-smod P1_P2_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;3328
                            end
                        end
                        else begin
                            $display(";A 3320");		//(= P1_P2_P3_Flush    0b0)) ;3320
                        end
                        if (((32'b00000000000000000000000000001111 - P1_P2_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 3330");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;3330
                            P1_P2_P3_State2 = 4'sb1000; $display(";A 3332");		//(= P1_P2_P3_State2    0b1000)) ;3332
                            P1_P2_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 3333");		//(= P1_P2_P3_InstQueueWr_Addr    0b00000)) ;3333
                        end
                        else begin
                            $display(";A 3331");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P1_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;3331
                            P1_P2_P3_State2 = 4'sb1001; $display(";A 3334");		//(= P1_P2_P3_State2    0b1001)) ;3334
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 3335");		//(= P1_P2_P3_State2    0b1000)) ;3335
                        if ((P1_P2_P3_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 3336");		//(= (bool-to-bv (bv-le P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;3336
                            P1_P2_P3_InstQueue[P1_P2_P3_InstQueueWr_Addr] = P1_P2_P3_InstQueue[P1_P2_P3_InstQueueRd_Addr]; $display(";A 3338");		//(= P1_P2_P3_InstQueue    ( P1_P2_P3_InstQueue P1_P2_P3_InstQueueRd_Addr ))) ;3338
                            P1_P2_P3_InstQueueRd_Addr = ((P1_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3339");		//(= P1_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3339
                            P1_P2_P3_InstQueueWr_Addr = ((P1_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 3340");		//(= P1_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P1_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;3340
                            P1_P2_P3_State2 = 4'sb1000; $display(";A 3341");		//(= P1_P2_P3_State2    0b1000)) ;3341
                        end
                        else begin
                            $display(";A 3337");		//(= (bool-to-bv (bv-le P1_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;3337
                            P1_P2_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 3342");		//(= P1_P2_P3_InstQueueRd_Addr    0b00000)) ;3342
                            P1_P2_P3_State2 = 4'sb1001; $display(";A 3343");		//(= P1_P2_P3_State2    0b1001)) ;3343
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 3344");		//(= P1_P2_P3_State2    0b1001)) ;3344
                        P1_P2_P3_rEIP <= #1 P1_P2_P3_PhyAddrPointer; $display(";A 3345");		//(= P1_P2_P3_rEIP    P1_P2_P3_PhyAddrPointer )) ;3345
                        P1_P2_P3_State2 = 4'sb0001; $display(";A 3346");		//(= P1_P2_P3_State2    0b0001)) ;3346
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:4940
    always @(posedge P1_P2_P3_RESET or posedge P1_P2_P3_CLOCK) begin
        if ((P1_P2_P3_RESET == 1'b1)) begin
            $display(";A 3347");		//(= (bv-comp P1_P2_P3_RESET  0b1)   0b1)) ;3347
            P1_P2_P3_ByteEnable <= #1 4'b0000; $display(";A 3349");		//(= P1_P2_P3_ByteEnable    0b0000)) ;3349
            P1_P2_P3_NonAligned <= #1 1'b0; $display(";A 3350");		//(= P1_P2_P3_NonAligned    0b0)) ;3350
        end
        else begin
            $display(";A 3348");		//(= (bv-comp P1_P2_P3_RESET  0b1)   0b0)) ;3348
            case (P1_P2_P3_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 3351");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000000)) ;3351
                        case ((P1_P2_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 3352");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;3352
                                    P1_P2_P3_ByteEnable <= #1 4'b1110; $display(";A 3353");		//(= P1_P2_P3_ByteEnable    0b1110)) ;3353
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 3354");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;3354
                                    P1_P2_P3_ByteEnable <= #1 4'b1101; $display(";A 3355");		//(= P1_P2_P3_ByteEnable    0b1101)) ;3355
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 3356");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;3356
                                    P1_P2_P3_ByteEnable <= #1 4'b1011; $display(";A 3357");		//(= P1_P2_P3_ByteEnable    0b1011)) ;3357
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 3358");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;3358
                                    P1_P2_P3_ByteEnable <= #1 4'b0111; $display(";A 3359");		//(= P1_P2_P3_ByteEnable    0b0111)) ;3359
                                end
                            default:
                                begin
                                    $display(";A 3360");		//(= (and (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;3360
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 3361");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000001)) ;3361
                        case ((P1_P2_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 3362");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;3362
                                    P1_P2_P3_ByteEnable <= #1 4'b1100; $display(";A 3363");		//(= P1_P2_P3_ByteEnable    0b1100)) ;3363
                                    P1_P2_P3_NonAligned <= #1 1'b0; $display(";A 3364");		//(= P1_P2_P3_NonAligned    0b0)) ;3364
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 3365");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;3365
                                    P1_P2_P3_ByteEnable <= #1 4'b1001; $display(";A 3366");		//(= P1_P2_P3_ByteEnable    0b1001)) ;3366
                                    P1_P2_P3_NonAligned <= #1 1'b0; $display(";A 3367");		//(= P1_P2_P3_NonAligned    0b0)) ;3367
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 3368");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;3368
                                    P1_P2_P3_ByteEnable <= #1 4'b0011; $display(";A 3369");		//(= P1_P2_P3_ByteEnable    0b0011)) ;3369
                                    P1_P2_P3_NonAligned <= #1 1'b0; $display(";A 3370");		//(= P1_P2_P3_NonAligned    0b0)) ;3370
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 3371");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;3371
                                    P1_P2_P3_ByteEnable <= #1 4'b0111; $display(";A 3372");		//(= P1_P2_P3_ByteEnable    0b0111)) ;3372
                                    P1_P2_P3_NonAligned <= #1 1'b1; $display(";A 3373");		//(= P1_P2_P3_NonAligned    0b1)) ;3373
                                end
                            default:
                                begin
                                    $display(";A 3374");		//(= (and (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;3374
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 3375");		//(= P1_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;3375
                        case ((P1_P2_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 3376");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;3376
                                    P1_P2_P3_ByteEnable <= #1 4'b0000; $display(";A 3377");		//(= P1_P2_P3_ByteEnable    0b0000)) ;3377
                                    P1_P2_P3_NonAligned <= #1 1'b0; $display(";A 3378");		//(= P1_P2_P3_NonAligned    0b0)) ;3378
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 3379");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;3379
                                    P1_P2_P3_ByteEnable <= #1 4'b0001; $display(";A 3380");		//(= P1_P2_P3_ByteEnable    0b0001)) ;3380
                                    P1_P2_P3_NonAligned <= #1 1'b1; $display(";A 3381");		//(= P1_P2_P3_NonAligned    0b1)) ;3381
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 3382");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;3382
                                    P1_P2_P3_NonAligned <= #1 1'b1; $display(";A 3383");		//(= P1_P2_P3_NonAligned    0b1)) ;3383
                                    P1_P2_P3_ByteEnable <= #1 4'b0011; $display(";A 3384");		//(= P1_P2_P3_ByteEnable    0b0011)) ;3384
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 3385");		//(= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;3385
                                    P1_P2_P3_NonAligned <= #1 1'b1; $display(";A 3386");		//(= P1_P2_P3_NonAligned    0b1)) ;3386
                                    P1_P2_P3_ByteEnable <= #1 4'b0111; $display(";A 3387");		//(= P1_P2_P3_ByteEnable    0b0111)) ;3387
                                end
                            default:
                                begin
                                    $display(";A 3388");		//(= (and (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P1_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;3388
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 3389");		//(= (and (/= P1_P2_P3_DataWidth  0b00000000000000000000000000000000) (/= P1_P2_P3_DataWidth  0b00000000000000000000000000000001) (/= P1_P2_P3_DataWidth  0b00000000000000000000000000000010))   true)) ;3389
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:5057
    always @(posedge P1_P3_reset or posedge P1_P3_clock) begin
        if ((P1_P3_reset == 1'b1)) begin
            P1_P3_MAR = 20'sb00000000000000000000; $display(";A 3392");		//(= P1_P3_MAR    0b00000000000000000000)) ;3392
            P1_P3_MBR = 32'sb00000000000000000000000000000000; $display(";A 3393");		//(= P1_P3_MBR    0b00000000000000000000000000000000)) ;3393
            P1_P3_IR = 32'sb00000000000000000000000000000000; $display(";A 3394");		//(= P1_P3_IR    0b00000000000000000000000000000000)) ;3394
            P1_P3_d = 32'sb00000000000000000000000000000000; $display(";A 3395");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3395
            P1_P3_r = 32'sb00000000000000000000000000000000; $display(";A 3396");		//(= P1_P3_r    0b00000000000000000000000000000000)) ;3396
            P1_P3_m = 32'sb00000000000000000000000000000000; $display(";A 3397");		//(= P1_P3_m    0b00000000000000000000000000000000)) ;3397
            P1_P3_s = 2'sb00; $display(";A 3398");		//(= P1_P3_s    0b00)) ;3398
            P1_P3_temp = 32'sb00000000000000000000000000000000; $display(";A 3399");		//(= P1_P3_temp    0b00000000000000000000000000000000)) ;3399
            P1_P3_mf = 2'sb00; $display(";A 3400");		//(= P1_P3_mf    0b00)) ;3400
            P1_P3_df = 3'sb000; $display(";A 3401");		//(= P1_P3_df    0b000)) ;3401
            P1_P3_ff = 4'sb0000; $display(";A 3402");		//(= P1_P3_ff    0b0000)) ;3402
            P1_P3_cf = 1'sb0; $display(";A 3403");		//(= P1_P3_cf    0b0)) ;3403
            P1_P3_tail = 20'sb00000000000000000000; $display(";A 3404");		//(= P1_P3_tail    0b00000000000000000000)) ;3404
            P1_P3_B = 1'b0; $display(";A 3405");		//(= P1_P3_B    0b0)) ;3405
            P1_P3_reg0 = 32'sb00000000000000000000000000000000; $display(";A 3406");		//(= P1_P3_reg0    0b00000000000000000000000000000000)) ;3406
            P1_P3_reg1 = 32'sb00000000000000000000000000000000; $display(";A 3407");		//(= P1_P3_reg1    0b00000000000000000000000000000000)) ;3407
            P1_P3_reg2 = 32'sb00000000000000000000000000000000; $display(";A 3408");		//(= P1_P3_reg2    0b00000000000000000000000000000000)) ;3408
            P1_P3_reg3 = 32'sb00000000000000000000000000000000; $display(";A 3409");		//(= P1_P3_reg3    0b00000000000000000000000000000000)) ;3409
            P1_P3_addr <= #1 20'sb00000000000000000000; $display(";A 3410");		//(= P1_P3_addr    0b00000000000000000000)) ;3410
            P1_P3_rd <= #1 1'b0; $display(";A 3411");		//(= P1_P3_rd    0b0)) ;3411
            P1_P3_wr <= #1 1'b0; $display(";A 3412");		//(= P1_P3_wr    0b0)) ;3412
            P1_P3_datao <= #1 32'sb00000000000000000000000000000000; $display(";A 3413");		//(= P1_P3_datao    0b00000000000000000000000000000000)) ;3413
            P1_P3_state = 1'sb0; $display(";A 3414");		//(= P1_P3_state    0b0)) ;3414
        end
        else begin
            P1_P3_rd <= #1 1'b0; $display(";A 3415");		//(= P1_P3_rd    0b0)) ;3415
            P1_P3_wr <= #1 1'b0; $display(";A 3416");		//(= P1_P3_wr    0b0)) ;3416
            case (P1_P3_state)
                1'b0 :
                    begin
                        $display(";A 3417");		//(= P1_P3_state    0b0)) ;3417
                        P1_P3_MAR = (P1_P3_reg3 % 32'b00000000000100000000000000000000); $display(";A 3418");		//(= P1_P3_MAR    (bv-smod P1_P3_reg3  0b00000000000100000000000000000000))) ;3418
                        P1_P3_addr <= #1 P1_P3_MAR; $display(";A 3419");		//(= P1_P3_addr    P1_P3_MAR )) ;3419
                        P1_P3_rd <= #1 1'b1; $display(";A 3420");		//(= P1_P3_rd    0b1)) ;3420
                        P1_P3_MBR = P1_P3_datai; $display(";A 3421");		//(= P1_P3_MBR    P1_P3_datai )) ;3421
                        P1_P3_IR = P1_P3_MBR; $display(";A 3422");		//(= P1_P3_IR    P1_P3_MBR )) ;3422
                        P1_P3_state = 1'sb1; $display(";A 3423");		//(= P1_P3_state    0b1)) ;3423
                    end
                1'b1 :
                    begin
                        $display(";A 3424");		//(= P1_P3_state    0b1)) ;3424
                        if ((P1_P3_IR < 32'sb00000000000000000000000000000000)) begin
                            $display(";A 3425");		//(= (bool-to-bv (bv-slt P1_P3_IR  0b00000000000000000000000000000000))   0b1)) ;3425
                            P1_P3_IR = (-P1_P3_IR); $display(";A 3427");		//(= P1_P3_IR    (bv-neg P1_P3_IR ))) ;3427
                        end
                        else begin
                            $display(";A 3426");		//(= (bool-to-bv (bv-slt P1_P3_IR  0b00000000000000000000000000000000))   0b0)) ;3426
                        end
                        P1_P3_mf = ((P1_P3_IR / 32'b00001000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 3428");		//(= P1_P3_mf    (bv-smod (bv-sdiv P1_P3_IR  0b00001000000000000000000000000000) 0b00000000000000000000000000000100))) ;3428
                        P1_P3_df = ((P1_P3_IR / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000000001000); $display(";A 3429");		//(= P1_P3_df    (bv-smod (bv-sdiv P1_P3_IR  0b00000001000000000000000000000000) 0b00000000000000000000000000001000))) ;3429
                        P1_P3_ff = ((P1_P3_IR / 32'b00000000000010000000000000000000) % 32'b00000000000000000000000000010000); $display(";A 3430");		//(= P1_P3_ff    (bv-smod (bv-sdiv P1_P3_IR  0b00000000000010000000000000000000) 0b00000000000000000000000000010000))) ;3430
                        P1_P3_cf = ((P1_P3_IR / 32'b00000000100000000000000000000000) % 32'b00000000000000000000000000000010); $display(";A 3431");		//(= P1_P3_cf    (bv-smod (bv-sdiv P1_P3_IR  0b00000000100000000000000000000000) 0b00000000000000000000000000000010))) ;3431
                        P1_P3_tail = (P1_P3_IR % 32'b00000000000100000000000000000000); $display(";A 3432");		//(= P1_P3_tail    (bv-smod P1_P3_IR  0b00000000000100000000000000000000))) ;3432
                        P1_P3_reg3 = ((P1_P3_reg3 % 32'b00100000000000000000000000000000) + 32'b00000000000000000000000000001000); $display(";A 3433");		//(= P1_P3_reg3    (bv-add (bv-smod P1_P3_reg3  0b00100000000000000000000000000000) 0b00000000000000000000000000001000))) ;3433
                        P1_P3_s = ((P1_P3_IR / 32'b00100000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 3434");		//(= P1_P3_s    (bv-smod (bv-sdiv P1_P3_IR  0b00100000000000000000000000000000) 0b00000000000000000000000000000100))) ;3434
                        case (P1_P3_s)
                            2'b00 :
                                begin
                                    $display(";A 3435");		//(= P1_P3_s    0b00)) ;3435
                                    P1_P3_r = P1_P3_reg0; $display(";A 3436");		//(= P1_P3_r    P1_P3_reg0 )) ;3436
                                end
                            2'b01 :
                                begin
                                    $display(";A 3437");		//(= P1_P3_s    0b01)) ;3437
                                    P1_P3_r = P1_P3_reg1; $display(";A 3438");		//(= P1_P3_r    P1_P3_reg1 )) ;3438
                                end
                            2'b10 :
                                begin
                                    $display(";A 3439");		//(= P1_P3_s    0b10)) ;3439
                                    P1_P3_r = P1_P3_reg2; $display(";A 3440");		//(= P1_P3_r    P1_P3_reg2 )) ;3440
                                end
                            2'b11 :
                                begin
                                    $display(";A 3441");		//(= P1_P3_s    0b11)) ;3441
                                    P1_P3_r = P1_P3_reg3; $display(";A 3442");		//(= P1_P3_r    P1_P3_reg3 )) ;3442
                                end
                        endcase
                        case (P1_P3_cf)
                            1'b1 :
                                begin
                                    $display(";A 3443");		//(= P1_P3_cf    0b1)) ;3443
                                    case (P1_P3_mf)
                                        2'b00 :
                                            begin
                                                $display(";A 3444");		//(= P1_P3_mf    0b00)) ;3444
                                                P1_P3_m = P1_P3_tail; $display(";A 3445");		//(= P1_P3_m    P1_P3_tail )) ;3445
                                            end
                                        2'b01 :
                                            begin
                                                $display(";A 3446");		//(= P1_P3_mf    0b01)) ;3446
                                                P1_P3_m = P1_P3_datai; $display(";A 3447");		//(= P1_P3_m    P1_P3_datai )) ;3447
                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3448");		//(= P1_P3_addr    P1_P3_tail )) ;3448
                                                P1_P3_rd <= #1 1'b1; $display(";A 3449");		//(= P1_P3_rd    0b1)) ;3449
                                            end
                                        2'b10 :
                                            begin
                                                $display(";A 3450");		//(= P1_P3_mf    0b10)) ;3450
                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3451");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3451
                                                P1_P3_rd <= #1 1'b1; $display(";A 3452");		//(= P1_P3_rd    0b1)) ;3452
                                                P1_P3_m = P1_P3_datai; $display(";A 3453");		//(= P1_P3_m    P1_P3_datai )) ;3453
                                            end
                                        2'b11 :
                                            begin
                                                $display(";A 3454");		//(= P1_P3_mf    0b11)) ;3454
                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3455");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3455
                                                P1_P3_rd <= #1 1'b1; $display(";A 3456");		//(= P1_P3_rd    0b1)) ;3456
                                                P1_P3_m = P1_P3_datai; $display(";A 3457");		//(= P1_P3_m    P1_P3_datai )) ;3457
                                            end
                                    endcase
                                    case (P1_P3_ff)
                                        4'b0000 :
                                            begin
                                                $display(";A 3458");		//(= P1_P3_ff    0b0000)) ;3458
                                                if ((P1_P3_r < P1_P3_m)) begin
                                                    $display(";A 3459");		//(= (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))   0b1)) ;3459
                                                    P1_P3_B = 1'b1; $display(";A 3461");		//(= P1_P3_B    0b1)) ;3461
                                                end
                                                else begin
                                                    $display(";A 3460");		//(= (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))   0b0)) ;3460
                                                    P1_P3_B = 1'b0; $display(";A 3462");		//(= P1_P3_B    0b0)) ;3462
                                                end
                                            end
                                        4'b0001 :
                                            begin
                                                $display(";A 3463");		//(= P1_P3_ff    0b0001)) ;3463
                                                if ((~(P1_P3_r < P1_P3_m))) begin
                                                    $display(";A 3464");		//(= (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )))   0b1)) ;3464
                                                    P1_P3_B = 1'b1; $display(";A 3466");		//(= P1_P3_B    0b1)) ;3466
                                                end
                                                else begin
                                                    $display(";A 3465");		//(= (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )))   0b0)) ;3465
                                                    P1_P3_B = 1'b0; $display(";A 3467");		//(= P1_P3_B    0b0)) ;3467
                                                end
                                            end
                                        4'b0010 :
                                            begin
                                                $display(";A 3468");		//(= P1_P3_ff    0b0010)) ;3468
                                                if ((P1_P3_r == P1_P3_m)) begin
                                                    $display(";A 3469");		//(= (bv-comp P1_P3_r  P1_P3_m )   0b1)) ;3469
                                                    P1_P3_B = 1'b1; $display(";A 3471");		//(= P1_P3_B    0b1)) ;3471
                                                end
                                                else begin
                                                    $display(";A 3470");		//(= (bv-comp P1_P3_r  P1_P3_m )   0b0)) ;3470
                                                    P1_P3_B = 1'b0; $display(";A 3472");		//(= P1_P3_B    0b0)) ;3472
                                                end
                                            end
                                        4'b0011 :
                                            begin
                                                $display(";A 3473");		//(= P1_P3_ff    0b0011)) ;3473
                                                if ((~(P1_P3_r == P1_P3_m))) begin
                                                    $display(";A 3474");		//(= (bv-not (bv-comp P1_P3_r  P1_P3_m ))   0b1)) ;3474
                                                    P1_P3_B = 1'b1; $display(";A 3476");		//(= P1_P3_B    0b1)) ;3476
                                                end
                                                else begin
                                                    $display(";A 3475");		//(= (bv-not (bv-comp P1_P3_r  P1_P3_m ))   0b0)) ;3475
                                                    P1_P3_B = 1'b0; $display(";A 3477");		//(= P1_P3_B    0b0)) ;3477
                                                end
                                            end
                                        4'b0100 :
                                            begin
                                                $display(";A 3478");		//(= P1_P3_ff    0b0100)) ;3478
                                                if ((~(P1_P3_r > P1_P3_m))) begin
                                                    $display(";A 3479");		//(= (bv-not (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m )))   0b1)) ;3479
                                                    P1_P3_B = 1'b1; $display(";A 3481");		//(= P1_P3_B    0b1)) ;3481
                                                end
                                                else begin
                                                    $display(";A 3480");		//(= (bv-not (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m )))   0b0)) ;3480
                                                    P1_P3_B = 1'b0; $display(";A 3482");		//(= P1_P3_B    0b0)) ;3482
                                                end
                                            end
                                        4'b0101 :
                                            begin
                                                $display(";A 3483");		//(= P1_P3_ff    0b0101)) ;3483
                                                if ((P1_P3_r > P1_P3_m)) begin
                                                    $display(";A 3484");		//(= (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m ))   0b1)) ;3484
                                                    P1_P3_B = 1'b1; $display(";A 3486");		//(= P1_P3_B    0b1)) ;3486
                                                end
                                                else begin
                                                    $display(";A 3485");		//(= (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m ))   0b0)) ;3485
                                                    P1_P3_B = 1'b0; $display(";A 3487");		//(= P1_P3_B    0b0)) ;3487
                                                end
                                            end
                                        4'b0110 :
                                            begin
                                                $display(";A 3488");		//(= P1_P3_ff    0b0110)) ;3488
                                                if ((P1_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 3489");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b1)) ;3489
                                                    P1_P3_r = (P1_P3_r - 32'b00000000000000000000000000000000); $display(";A 3491");		//(= P1_P3_r    (bv-sub P1_P3_r  0b00000000000000000000000000000000))) ;3491
                                                end
                                                else begin
                                                    $display(";A 3490");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b0)) ;3490
                                                end
                                                if ((P1_P3_r < P1_P3_m)) begin
                                                    $display(";A 3492");		//(= (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))   0b1)) ;3492
                                                    P1_P3_B = 1'b1; $display(";A 3494");		//(= P1_P3_B    0b1)) ;3494
                                                end
                                                else begin
                                                    $display(";A 3493");		//(= (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))   0b0)) ;3493
                                                    P1_P3_B = 1'b0; $display(";A 3495");		//(= P1_P3_B    0b0)) ;3495
                                                end
                                            end
                                        4'b0111 :
                                            begin
                                                $display(";A 3496");		//(= P1_P3_ff    0b0111)) ;3496
                                                if ((P1_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 3497");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b1)) ;3497
                                                    P1_P3_r = (P1_P3_r - 32'b00000000000000000000000000000000); $display(";A 3499");		//(= P1_P3_r    (bv-sub P1_P3_r  0b00000000000000000000000000000000))) ;3499
                                                end
                                                else begin
                                                    $display(";A 3498");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b0)) ;3498
                                                end
                                                if ((~(P1_P3_r < P1_P3_m))) begin
                                                    $display(";A 3500");		//(= (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )))   0b1)) ;3500
                                                    P1_P3_B = 1'b1; $display(";A 3502");		//(= P1_P3_B    0b1)) ;3502
                                                end
                                                else begin
                                                    $display(";A 3501");		//(= (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )))   0b0)) ;3501
                                                    P1_P3_B = 1'b0; $display(";A 3503");		//(= P1_P3_B    0b0)) ;3503
                                                end
                                            end
                                        4'b1000 :
                                            begin
                                                $display(";A 3504");		//(= P1_P3_ff    0b1000)) ;3504
                                                if (((P1_P3_r < P1_P3_m) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3505");		//(= (bv-or (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b1)) ;3505
                                                    P1_P3_B = 1'b1; $display(";A 3507");		//(= P1_P3_B    0b1)) ;3507
                                                end
                                                else begin
                                                    $display(";A 3506");		//(= (bv-or (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b0)) ;3506
                                                    P1_P3_B = 1'b0; $display(";A 3508");		//(= P1_P3_B    0b0)) ;3508
                                                end
                                            end
                                        4'b1001 :
                                            begin
                                                $display(";A 3509");		//(= P1_P3_ff    0b1001)) ;3509
                                                if (((~(P1_P3_r < P1_P3_m)) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3510");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))) (bv-comp P1_P3_B  0b1))   0b1)) ;3510
                                                    P1_P3_B = 1'b1; $display(";A 3512");		//(= P1_P3_B    0b1)) ;3512
                                                end
                                                else begin
                                                    $display(";A 3511");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))) (bv-comp P1_P3_B  0b1))   0b0)) ;3511
                                                    P1_P3_B = 1'b0; $display(";A 3513");		//(= P1_P3_B    0b0)) ;3513
                                                end
                                            end
                                        4'b1010 :
                                            begin
                                                $display(";A 3514");		//(= P1_P3_ff    0b1010)) ;3514
                                                if (((P1_P3_r == P1_P3_m) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3515");		//(= (bv-or (bv-comp P1_P3_r  P1_P3_m ) (bv-comp P1_P3_B  0b1))   0b1)) ;3515
                                                    P1_P3_B = 1'b1; $display(";A 3517");		//(= P1_P3_B    0b1)) ;3517
                                                end
                                                else begin
                                                    $display(";A 3516");		//(= (bv-or (bv-comp P1_P3_r  P1_P3_m ) (bv-comp P1_P3_B  0b1))   0b0)) ;3516
                                                    P1_P3_B = 1'b0; $display(";A 3518");		//(= P1_P3_B    0b0)) ;3518
                                                end
                                            end
                                        4'b1011 :
                                            begin
                                                $display(";A 3519");		//(= P1_P3_ff    0b1011)) ;3519
                                                if (((~(P1_P3_r == P1_P3_m)) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3520");		//(= (bv-or (bv-not (bv-comp P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b1)) ;3520
                                                    P1_P3_B = 1'b1; $display(";A 3522");		//(= P1_P3_B    0b1)) ;3522
                                                end
                                                else begin
                                                    $display(";A 3521");		//(= (bv-or (bv-not (bv-comp P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b0)) ;3521
                                                    P1_P3_B = 1'b0; $display(";A 3523");		//(= P1_P3_B    0b0)) ;3523
                                                end
                                            end
                                        4'b1100 :
                                            begin
                                                $display(";A 3524");		//(= P1_P3_ff    0b1100)) ;3524
                                                if (((~(P1_P3_r > P1_P3_m)) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3525");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m ))) (bv-comp P1_P3_B  0b1))   0b1)) ;3525
                                                    P1_P3_B = 1'b1; $display(";A 3527");		//(= P1_P3_B    0b1)) ;3527
                                                end
                                                else begin
                                                    $display(";A 3526");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m ))) (bv-comp P1_P3_B  0b1))   0b0)) ;3526
                                                    P1_P3_B = 1'b0; $display(";A 3528");		//(= P1_P3_B    0b0)) ;3528
                                                end
                                            end
                                        4'b1101 :
                                            begin
                                                $display(";A 3529");		//(= P1_P3_ff    0b1101)) ;3529
                                                if (((P1_P3_r > P1_P3_m) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3530");		//(= (bv-or (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b1)) ;3530
                                                    P1_P3_B = 1'b1; $display(";A 3532");		//(= P1_P3_B    0b1)) ;3532
                                                end
                                                else begin
                                                    $display(";A 3531");		//(= (bv-or (bool-to-bv (bv-sgt P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b0)) ;3531
                                                    P1_P3_B = 1'b0; $display(";A 3533");		//(= P1_P3_B    0b0)) ;3533
                                                end
                                            end
                                        4'b1110 :
                                            begin
                                                $display(";A 3534");		//(= P1_P3_ff    0b1110)) ;3534
                                                if ((P1_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 3535");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b1)) ;3535
                                                    P1_P3_r = (P1_P3_r - 32'b00000000000000000000000000000000); $display(";A 3537");		//(= P1_P3_r    (bv-sub P1_P3_r  0b00000000000000000000000000000000))) ;3537
                                                end
                                                else begin
                                                    $display(";A 3536");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b0)) ;3536
                                                end
                                                if (((P1_P3_r < P1_P3_m) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3538");		//(= (bv-or (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b1)) ;3538
                                                    P1_P3_B = 1'b1; $display(";A 3540");		//(= P1_P3_B    0b1)) ;3540
                                                end
                                                else begin
                                                    $display(";A 3539");		//(= (bv-or (bool-to-bv (bv-slt P1_P3_r  P1_P3_m )) (bv-comp P1_P3_B  0b1))   0b0)) ;3539
                                                    P1_P3_B = 1'b0; $display(";A 3541");		//(= P1_P3_B    0b0)) ;3541
                                                end
                                            end
                                        4'b1111 :
                                            begin
                                                $display(";A 3542");		//(= P1_P3_ff    0b1111)) ;3542
                                                if ((P1_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 3543");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b1)) ;3543
                                                    P1_P3_r = (P1_P3_r - 32'b00000000000000000000000000000000); $display(";A 3545");		//(= P1_P3_r    (bv-sub P1_P3_r  0b00000000000000000000000000000000))) ;3545
                                                end
                                                else begin
                                                    $display(";A 3544");		//(= (bool-to-bv (bv-gt P1_P3_r  0b11111111111111111111111111111111))   0b0)) ;3544
                                                end
                                                if (((~(P1_P3_r < P1_P3_m)) | (P1_P3_B == 1'b1))) begin
                                                    $display(";A 3546");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))) (bv-comp P1_P3_B  0b1))   0b1)) ;3546
                                                    P1_P3_B = 1'b1; $display(";A 3548");		//(= P1_P3_B    0b1)) ;3548
                                                end
                                                else begin
                                                    $display(";A 3547");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P3_r  P1_P3_m ))) (bv-comp P1_P3_B  0b1))   0b0)) ;3547
                                                    P1_P3_B = 1'b0; $display(";A 3549");		//(= P1_P3_B    0b0)) ;3549
                                                end
                                            end
                                    endcase
                                end
                            1'b0 :
                                begin
                                    $display(";A 3550");		//(= P1_P3_cf    0b0)) ;3550
                                    if ((~(P1_P3_df == 32'b00000000000000000000000000000111))) begin
                                        $display(";A 3551");		//(= (bv-not (bv-comp P1_P3_df  0b00000000000000000000000000000111))   0b1)) ;3551
                                        if ((P1_P3_df == 32'b00000000000000000000000000000101)) begin
                                            $display(";A 3553");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000101)   0b1)) ;3553
                                            if (((~P1_P3_B) == 1'b1)) begin
                                                $display(";A 3555");		//(= (bv-comp (bv-not P1_P3_B ) 0b1)   0b1)) ;3555
                                                P1_P3_d = 32'sb00000000000000000000000000000011; $display(";A 3557");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3557
                                            end
                                            else begin
                                                $display(";A 3556");		//(= (bv-comp (bv-not P1_P3_B ) 0b1)   0b0)) ;3556
                                            end
                                        end
                                        else begin
                                            $display(";A 3554");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000101)   0b0)) ;3554
                                            if ((P1_P3_df == 32'b00000000000000000000000000000100)) begin
                                                $display(";A 3558");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000100)   0b1)) ;3558
                                                if ((P1_P3_B == 1'b1)) begin
                                                    $display(";A 3560");		//(= (bv-comp P1_P3_B  0b1)   0b1)) ;3560
                                                    P1_P3_d = 32'sb00000000000000000000000000000011; $display(";A 3562");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3562
                                                end
                                                else begin
                                                    $display(";A 3561");		//(= (bv-comp P1_P3_B  0b1)   0b0)) ;3561
                                                end
                                            end
                                            else begin
                                                $display(";A 3559");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000100)   0b0)) ;3559
                                                if ((P1_P3_df == 32'b00000000000000000000000000000011)) begin
                                                    $display(";A 3563");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000011)   0b1)) ;3563
                                                    P1_P3_d = 32'sb00000000000000000000000000000011; $display(";A 3565");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3565
                                                end
                                                else begin
                                                    $display(";A 3564");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000011)   0b0)) ;3564
                                                    if ((P1_P3_df == 32'b00000000000000000000000000000010)) begin
                                                        $display(";A 3566");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000010)   0b1)) ;3566
                                                        P1_P3_d = 32'sb00000000000000000000000000000010; $display(";A 3568");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3568
                                                    end
                                                    else begin
                                                        $display(";A 3567");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000010)   0b0)) ;3567
                                                        if ((P1_P3_df == 32'b00000000000000000000000000000001)) begin
                                                            $display(";A 3569");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000001)   0b1)) ;3569
                                                            P1_P3_d = 32'sb00000000000000000000000000000001; $display(";A 3571");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3571
                                                        end
                                                        else begin
                                                            $display(";A 3570");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000001)   0b0)) ;3570
                                                            if ((P1_P3_df == 32'b00000000000000000000000000000000)) begin
                                                                $display(";A 3572");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000000)   0b1)) ;3572
                                                                P1_P3_d = 32'sb00000000000000000000000000000000; $display(";A 3574");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3574
                                                            end
                                                            else begin
                                                                $display(";A 3573");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000000)   0b0)) ;3573
                                                            end
                                                        end
                                                    end
                                                end
                                            end
                                        end
                                        case (P1_P3_ff)
                                            4'b0000 :
                                                begin
                                                    $display(";A 3575");		//(= P1_P3_ff    0b0000)) ;3575
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3576");		//(= P1_P3_mf    0b00)) ;3576
                                                                P1_P3_m = P1_P3_tail; $display(";A 3577");		//(= P1_P3_m    P1_P3_tail )) ;3577
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3578");		//(= P1_P3_mf    0b01)) ;3578
                                                                P1_P3_m = P1_P3_datai; $display(";A 3579");		//(= P1_P3_m    P1_P3_datai )) ;3579
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3580");		//(= P1_P3_addr    P1_P3_tail )) ;3580
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3581");		//(= P1_P3_rd    0b1)) ;3581
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3582");		//(= P1_P3_mf    0b10)) ;3582
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3583");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3583
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3584");		//(= P1_P3_rd    0b1)) ;3584
                                                                P1_P3_m = P1_P3_datai; $display(";A 3585");		//(= P1_P3_m    P1_P3_datai )) ;3585
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3586");		//(= P1_P3_mf    0b11)) ;3586
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3587");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3587
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3588");		//(= P1_P3_rd    0b1)) ;3588
                                                                P1_P3_m = P1_P3_datai; $display(";A 3589");		//(= P1_P3_m    P1_P3_datai )) ;3589
                                                            end
                                                    endcase
                                                    P1_P3_t = 32'sb00000000000000000000000000000000; $display(";A 3590");		//(= P1_P3_t    0b00000000000000000000000000000000)) ;3590
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3591");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3591
                                                                P1_P3_reg0 = (P1_P3_t - P1_P3_m); $display(";A 3592");		//(= P1_P3_reg0    (bv-sub P1_P3_t  P1_P3_m ))) ;3592
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3593");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3593
                                                                P1_P3_reg1 = (P1_P3_t - P1_P3_m); $display(";A 3594");		//(= P1_P3_reg1    (bv-sub P1_P3_t  P1_P3_m ))) ;3594
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3595");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3595
                                                                P1_P3_reg2 = (P1_P3_t - P1_P3_m); $display(";A 3596");		//(= P1_P3_reg2    (bv-sub P1_P3_t  P1_P3_m ))) ;3596
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3597");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3597
                                                                P1_P3_reg3 = (P1_P3_t - P1_P3_m); $display(";A 3598");		//(= P1_P3_reg3    (bv-sub P1_P3_t  P1_P3_m ))) ;3598
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3599");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3599
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0001 :
                                                begin
                                                    $display(";A 3600");		//(= P1_P3_ff    0b0001)) ;3600
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3601");		//(= P1_P3_mf    0b00)) ;3601
                                                                P1_P3_m = P1_P3_tail; $display(";A 3602");		//(= P1_P3_m    P1_P3_tail )) ;3602
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3603");		//(= P1_P3_mf    0b01)) ;3603
                                                                P1_P3_m = P1_P3_datai; $display(";A 3604");		//(= P1_P3_m    P1_P3_datai )) ;3604
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3605");		//(= P1_P3_addr    P1_P3_tail )) ;3605
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3606");		//(= P1_P3_rd    0b1)) ;3606
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3607");		//(= P1_P3_mf    0b10)) ;3607
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3608");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3608
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3609");		//(= P1_P3_rd    0b1)) ;3609
                                                                P1_P3_m = P1_P3_datai; $display(";A 3610");		//(= P1_P3_m    P1_P3_datai )) ;3610
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3611");		//(= P1_P3_mf    0b11)) ;3611
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3612");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3612
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3613");		//(= P1_P3_rd    0b1)) ;3613
                                                                P1_P3_m = P1_P3_datai; $display(";A 3614");		//(= P1_P3_m    P1_P3_datai )) ;3614
                                                            end
                                                    endcase
                                                    P1_P3_reg2 = P1_P3_reg3; $display(";A 3615");		//(= P1_P3_reg2    P1_P3_reg3 )) ;3615
                                                    P1_P3_reg3 = P1_P3_m; $display(";A 3616");		//(= P1_P3_reg3    P1_P3_m )) ;3616
                                                end
                                            4'b0010 :
                                                begin
                                                    $display(";A 3617");		//(= P1_P3_ff    0b0010)) ;3617
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3618");		//(= P1_P3_mf    0b00)) ;3618
                                                                P1_P3_m = P1_P3_tail; $display(";A 3619");		//(= P1_P3_m    P1_P3_tail )) ;3619
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3620");		//(= P1_P3_mf    0b01)) ;3620
                                                                P1_P3_m = P1_P3_datai; $display(";A 3621");		//(= P1_P3_m    P1_P3_datai )) ;3621
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3622");		//(= P1_P3_addr    P1_P3_tail )) ;3622
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3623");		//(= P1_P3_rd    0b1)) ;3623
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3624");		//(= P1_P3_mf    0b10)) ;3624
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3625");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3625
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3626");		//(= P1_P3_rd    0b1)) ;3626
                                                                P1_P3_m = P1_P3_datai; $display(";A 3627");		//(= P1_P3_m    P1_P3_datai )) ;3627
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3628");		//(= P1_P3_mf    0b11)) ;3628
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3629");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3629
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3630");		//(= P1_P3_rd    0b1)) ;3630
                                                                P1_P3_m = P1_P3_datai; $display(";A 3631");		//(= P1_P3_m    P1_P3_datai )) ;3631
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3632");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3632
                                                                P1_P3_reg0 = P1_P3_m; $display(";A 3633");		//(= P1_P3_reg0    P1_P3_m )) ;3633
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3634");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3634
                                                                P1_P3_reg1 = P1_P3_m; $display(";A 3635");		//(= P1_P3_reg1    P1_P3_m )) ;3635
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3636");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3636
                                                                P1_P3_reg2 = P1_P3_m; $display(";A 3637");		//(= P1_P3_reg2    P1_P3_m )) ;3637
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3638");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3638
                                                                P1_P3_reg3 = P1_P3_m; $display(";A 3639");		//(= P1_P3_reg3    P1_P3_m )) ;3639
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3640");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3640
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0011 :
                                                begin
                                                    $display(";A 3641");		//(= P1_P3_ff    0b0011)) ;3641
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3642");		//(= P1_P3_mf    0b00)) ;3642
                                                                P1_P3_m = P1_P3_tail; $display(";A 3643");		//(= P1_P3_m    P1_P3_tail )) ;3643
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3644");		//(= P1_P3_mf    0b01)) ;3644
                                                                P1_P3_m = P1_P3_datai; $display(";A 3645");		//(= P1_P3_m    P1_P3_datai )) ;3645
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3646");		//(= P1_P3_addr    P1_P3_tail )) ;3646
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3647");		//(= P1_P3_rd    0b1)) ;3647
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3648");		//(= P1_P3_mf    0b10)) ;3648
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3649");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3649
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3650");		//(= P1_P3_rd    0b1)) ;3650
                                                                P1_P3_m = P1_P3_datai; $display(";A 3651");		//(= P1_P3_m    P1_P3_datai )) ;3651
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3652");		//(= P1_P3_mf    0b11)) ;3652
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3653");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3653
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3654");		//(= P1_P3_rd    0b1)) ;3654
                                                                P1_P3_m = P1_P3_datai; $display(";A 3655");		//(= P1_P3_m    P1_P3_datai )) ;3655
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3656");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3656
                                                                P1_P3_reg0 = P1_P3_m; $display(";A 3657");		//(= P1_P3_reg0    P1_P3_m )) ;3657
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3658");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3658
                                                                P1_P3_reg1 = P1_P3_m; $display(";A 3659");		//(= P1_P3_reg1    P1_P3_m )) ;3659
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3660");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3660
                                                                P1_P3_reg2 = P1_P3_m; $display(";A 3661");		//(= P1_P3_reg2    P1_P3_m )) ;3661
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3662");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3662
                                                                P1_P3_reg3 = P1_P3_m; $display(";A 3663");		//(= P1_P3_reg3    P1_P3_m )) ;3663
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3664");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3664
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0100 :
                                                begin
                                                    $display(";A 3665");		//(= P1_P3_ff    0b0100)) ;3665
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3666");		//(= P1_P3_mf    0b00)) ;3666
                                                                P1_P3_m = P1_P3_tail; $display(";A 3667");		//(= P1_P3_m    P1_P3_tail )) ;3667
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3668");		//(= P1_P3_mf    0b01)) ;3668
                                                                P1_P3_m = P1_P3_datai; $display(";A 3669");		//(= P1_P3_m    P1_P3_datai )) ;3669
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3670");		//(= P1_P3_addr    P1_P3_tail )) ;3670
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3671");		//(= P1_P3_rd    0b1)) ;3671
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3672");		//(= P1_P3_mf    0b10)) ;3672
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3673");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3673
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3674");		//(= P1_P3_rd    0b1)) ;3674
                                                                P1_P3_m = P1_P3_datai; $display(";A 3675");		//(= P1_P3_m    P1_P3_datai )) ;3675
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3676");		//(= P1_P3_mf    0b11)) ;3676
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3677");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3677
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3678");		//(= P1_P3_rd    0b1)) ;3678
                                                                P1_P3_m = P1_P3_datai; $display(";A 3679");		//(= P1_P3_m    P1_P3_datai )) ;3679
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3680");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3680
                                                                P1_P3_reg0 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3681");		//(= P1_P3_reg0    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3681
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3682");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3682
                                                                P1_P3_reg1 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3683");		//(= P1_P3_reg1    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3683
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3684");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3684
                                                                P1_P3_reg2 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3685");		//(= P1_P3_reg2    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3685
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3686");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3686
                                                                P1_P3_reg3 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3687");		//(= P1_P3_reg3    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3687
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3688");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3688
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0101 :
                                                begin
                                                    $display(";A 3689");		//(= P1_P3_ff    0b0101)) ;3689
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3690");		//(= P1_P3_mf    0b00)) ;3690
                                                                P1_P3_m = P1_P3_tail; $display(";A 3691");		//(= P1_P3_m    P1_P3_tail )) ;3691
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3692");		//(= P1_P3_mf    0b01)) ;3692
                                                                P1_P3_m = P1_P3_datai; $display(";A 3693");		//(= P1_P3_m    P1_P3_datai )) ;3693
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3694");		//(= P1_P3_addr    P1_P3_tail )) ;3694
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3695");		//(= P1_P3_rd    0b1)) ;3695
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3696");		//(= P1_P3_mf    0b10)) ;3696
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3697");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3697
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3698");		//(= P1_P3_rd    0b1)) ;3698
                                                                P1_P3_m = P1_P3_datai; $display(";A 3699");		//(= P1_P3_m    P1_P3_datai )) ;3699
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3700");		//(= P1_P3_mf    0b11)) ;3700
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3701");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3701
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3702");		//(= P1_P3_rd    0b1)) ;3702
                                                                P1_P3_m = P1_P3_datai; $display(";A 3703");		//(= P1_P3_m    P1_P3_datai )) ;3703
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3704");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3704
                                                                P1_P3_reg0 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3705");		//(= P1_P3_reg0    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3705
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3706");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3706
                                                                P1_P3_reg1 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3707");		//(= P1_P3_reg1    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3707
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3708");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3708
                                                                P1_P3_reg2 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3709");		//(= P1_P3_reg2    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3709
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3710");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3710
                                                                P1_P3_reg3 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3711");		//(= P1_P3_reg3    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3711
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3712");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3712
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0110 :
                                                begin
                                                    $display(";A 3713");		//(= P1_P3_ff    0b0110)) ;3713
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3714");		//(= P1_P3_mf    0b00)) ;3714
                                                                P1_P3_m = P1_P3_tail; $display(";A 3715");		//(= P1_P3_m    P1_P3_tail )) ;3715
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3716");		//(= P1_P3_mf    0b01)) ;3716
                                                                P1_P3_m = P1_P3_datai; $display(";A 3717");		//(= P1_P3_m    P1_P3_datai )) ;3717
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3718");		//(= P1_P3_addr    P1_P3_tail )) ;3718
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3719");		//(= P1_P3_rd    0b1)) ;3719
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3720");		//(= P1_P3_mf    0b10)) ;3720
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3721");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3721
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3722");		//(= P1_P3_rd    0b1)) ;3722
                                                                P1_P3_m = P1_P3_datai; $display(";A 3723");		//(= P1_P3_m    P1_P3_datai )) ;3723
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3724");		//(= P1_P3_mf    0b11)) ;3724
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3725");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3725
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3726");		//(= P1_P3_rd    0b1)) ;3726
                                                                P1_P3_m = P1_P3_datai; $display(";A 3727");		//(= P1_P3_m    P1_P3_datai )) ;3727
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3728");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3728
                                                                P1_P3_reg0 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3729");		//(= P1_P3_reg0    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3729
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3730");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3730
                                                                P1_P3_reg1 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3731");		//(= P1_P3_reg1    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3731
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3732");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3732
                                                                P1_P3_reg2 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3733");		//(= P1_P3_reg2    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3733
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3734");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3734
                                                                P1_P3_reg3 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3735");		//(= P1_P3_reg3    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3735
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3736");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3736
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0111 :
                                                begin
                                                    $display(";A 3737");		//(= P1_P3_ff    0b0111)) ;3737
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3738");		//(= P1_P3_mf    0b00)) ;3738
                                                                P1_P3_m = P1_P3_tail; $display(";A 3739");		//(= P1_P3_m    P1_P3_tail )) ;3739
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3740");		//(= P1_P3_mf    0b01)) ;3740
                                                                P1_P3_m = P1_P3_datai; $display(";A 3741");		//(= P1_P3_m    P1_P3_datai )) ;3741
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3742");		//(= P1_P3_addr    P1_P3_tail )) ;3742
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3743");		//(= P1_P3_rd    0b1)) ;3743
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3744");		//(= P1_P3_mf    0b10)) ;3744
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3745");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3745
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3746");		//(= P1_P3_rd    0b1)) ;3746
                                                                P1_P3_m = P1_P3_datai; $display(";A 3747");		//(= P1_P3_m    P1_P3_datai )) ;3747
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3748");		//(= P1_P3_mf    0b11)) ;3748
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3749");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3749
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3750");		//(= P1_P3_rd    0b1)) ;3750
                                                                P1_P3_m = P1_P3_datai; $display(";A 3751");		//(= P1_P3_m    P1_P3_datai )) ;3751
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3752");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3752
                                                                P1_P3_reg0 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3753");		//(= P1_P3_reg0    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3753
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3754");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3754
                                                                P1_P3_reg1 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3755");		//(= P1_P3_reg1    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3755
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3756");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3756
                                                                P1_P3_reg2 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3757");		//(= P1_P3_reg2    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3757
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3758");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3758
                                                                P1_P3_reg3 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3759");		//(= P1_P3_reg3    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3759
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3760");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3760
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1000 :
                                                begin
                                                    $display(";A 3761");		//(= P1_P3_ff    0b1000)) ;3761
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3762");		//(= P1_P3_mf    0b00)) ;3762
                                                                P1_P3_m = P1_P3_tail; $display(";A 3763");		//(= P1_P3_m    P1_P3_tail )) ;3763
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3764");		//(= P1_P3_mf    0b01)) ;3764
                                                                P1_P3_m = P1_P3_datai; $display(";A 3765");		//(= P1_P3_m    P1_P3_datai )) ;3765
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3766");		//(= P1_P3_addr    P1_P3_tail )) ;3766
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3767");		//(= P1_P3_rd    0b1)) ;3767
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3768");		//(= P1_P3_mf    0b10)) ;3768
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3769");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3769
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3770");		//(= P1_P3_rd    0b1)) ;3770
                                                                P1_P3_m = P1_P3_datai; $display(";A 3771");		//(= P1_P3_m    P1_P3_datai )) ;3771
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3772");		//(= P1_P3_mf    0b11)) ;3772
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3773");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3773
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3774");		//(= P1_P3_rd    0b1)) ;3774
                                                                P1_P3_m = P1_P3_datai; $display(";A 3775");		//(= P1_P3_m    P1_P3_datai )) ;3775
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3776");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3776
                                                                P1_P3_reg0 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3777");		//(= P1_P3_reg0    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3777
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3778");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3778
                                                                P1_P3_reg1 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3779");		//(= P1_P3_reg1    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3779
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3780");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3780
                                                                P1_P3_reg2 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3781");		//(= P1_P3_reg2    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3781
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3782");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3782
                                                                P1_P3_reg3 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3783");		//(= P1_P3_reg3    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3783
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3784");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3784
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1001 :
                                                begin
                                                    $display(";A 3785");		//(= P1_P3_ff    0b1001)) ;3785
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3786");		//(= P1_P3_mf    0b00)) ;3786
                                                                P1_P3_m = P1_P3_tail; $display(";A 3787");		//(= P1_P3_m    P1_P3_tail )) ;3787
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3788");		//(= P1_P3_mf    0b01)) ;3788
                                                                P1_P3_m = P1_P3_datai; $display(";A 3789");		//(= P1_P3_m    P1_P3_datai )) ;3789
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3790");		//(= P1_P3_addr    P1_P3_tail )) ;3790
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3791");		//(= P1_P3_rd    0b1)) ;3791
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3792");		//(= P1_P3_mf    0b10)) ;3792
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3793");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3793
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3794");		//(= P1_P3_rd    0b1)) ;3794
                                                                P1_P3_m = P1_P3_datai; $display(";A 3795");		//(= P1_P3_m    P1_P3_datai )) ;3795
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3796");		//(= P1_P3_mf    0b11)) ;3796
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3797");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3797
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3798");		//(= P1_P3_rd    0b1)) ;3798
                                                                P1_P3_m = P1_P3_datai; $display(";A 3799");		//(= P1_P3_m    P1_P3_datai )) ;3799
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3800");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3800
                                                                P1_P3_reg0 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3801");		//(= P1_P3_reg0    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3801
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3802");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3802
                                                                P1_P3_reg1 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3803");		//(= P1_P3_reg1    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3803
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3804");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3804
                                                                P1_P3_reg2 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3805");		//(= P1_P3_reg2    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3805
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3806");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3806
                                                                P1_P3_reg3 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3807");		//(= P1_P3_reg3    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3807
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3808");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3808
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1010 :
                                                begin
                                                    $display(";A 3809");		//(= P1_P3_ff    0b1010)) ;3809
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3810");		//(= P1_P3_mf    0b00)) ;3810
                                                                P1_P3_m = P1_P3_tail; $display(";A 3811");		//(= P1_P3_m    P1_P3_tail )) ;3811
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3812");		//(= P1_P3_mf    0b01)) ;3812
                                                                P1_P3_m = P1_P3_datai; $display(";A 3813");		//(= P1_P3_m    P1_P3_datai )) ;3813
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3814");		//(= P1_P3_addr    P1_P3_tail )) ;3814
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3815");		//(= P1_P3_rd    0b1)) ;3815
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3816");		//(= P1_P3_mf    0b10)) ;3816
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3817");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3817
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3818");		//(= P1_P3_rd    0b1)) ;3818
                                                                P1_P3_m = P1_P3_datai; $display(";A 3819");		//(= P1_P3_m    P1_P3_datai )) ;3819
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3820");		//(= P1_P3_mf    0b11)) ;3820
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3821");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3821
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3822");		//(= P1_P3_rd    0b1)) ;3822
                                                                P1_P3_m = P1_P3_datai; $display(";A 3823");		//(= P1_P3_m    P1_P3_datai )) ;3823
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3824");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3824
                                                                P1_P3_reg0 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3825");		//(= P1_P3_reg0    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3825
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3826");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3826
                                                                P1_P3_reg1 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3827");		//(= P1_P3_reg1    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3827
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3828");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3828
                                                                P1_P3_reg2 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3829");		//(= P1_P3_reg2    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3829
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3830");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3830
                                                                P1_P3_reg3 = ((P1_P3_r + P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3831");		//(= P1_P3_reg3    (bv-smod (bv-add P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3831
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3832");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3832
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1011 :
                                                begin
                                                    $display(";A 3833");		//(= P1_P3_ff    0b1011)) ;3833
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3834");		//(= P1_P3_mf    0b00)) ;3834
                                                                P1_P3_m = P1_P3_tail; $display(";A 3835");		//(= P1_P3_m    P1_P3_tail )) ;3835
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3836");		//(= P1_P3_mf    0b01)) ;3836
                                                                P1_P3_m = P1_P3_datai; $display(";A 3837");		//(= P1_P3_m    P1_P3_datai )) ;3837
                                                                P1_P3_addr <= #1 P1_P3_tail; $display(";A 3838");		//(= P1_P3_addr    P1_P3_tail )) ;3838
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3839");		//(= P1_P3_rd    0b1)) ;3839
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3840");		//(= P1_P3_mf    0b10)) ;3840
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 3841");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg1 ) 0b00000000000100000000000000000000))) ;3841
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3842");		//(= P1_P3_rd    0b1)) ;3842
                                                                P1_P3_m = P1_P3_datai; $display(";A 3843");		//(= P1_P3_m    P1_P3_datai )) ;3843
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3844");		//(= P1_P3_mf    0b11)) ;3844
                                                                P1_P3_addr <= #1 ((P1_P3_tail + P1_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 3845");		//(= P1_P3_addr    (bv-smod (bv-add P1_P3_tail  P1_P3_reg2 ) 0b00000000000100000000000000000000))) ;3845
                                                                P1_P3_rd <= #1 1'b1; $display(";A 3846");		//(= P1_P3_rd    0b1)) ;3846
                                                                P1_P3_m = P1_P3_datai; $display(";A 3847");		//(= P1_P3_m    P1_P3_datai )) ;3847
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3848");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3848
                                                                P1_P3_reg0 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3849");		//(= P1_P3_reg0    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3849
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3850");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3850
                                                                P1_P3_reg1 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3851");		//(= P1_P3_reg1    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3851
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3852");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3852
                                                                P1_P3_reg2 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3853");		//(= P1_P3_reg2    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3853
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3854");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3854
                                                                P1_P3_reg3 = ((P1_P3_r - P1_P3_m) % 32'b00000000000000000000000000000000); $display(";A 3855");		//(= P1_P3_reg3    (bv-smod (bv-sub P1_P3_r  P1_P3_m ) 0b00000000000000000000000000000000))) ;3855
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3856");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3856
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1100 :
                                                begin
                                                    $display(";A 3857");		//(= P1_P3_ff    0b1100)) ;3857
                                                    case (P1_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 3858");		//(= P1_P3_mf    0b00)) ;3858
                                                                P1_P3_t = (P1_P3_r / 32'sb00000000000000000000000000000010); $display(";A 3859");		//(= P1_P3_t    (bv-sdiv P1_P3_r  0b00000000000000000000000000000010))) ;3859
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 3860");		//(= P1_P3_mf    0b01)) ;3860
                                                                P1_P3_t = (P1_P3_r / 32'sb00000000000000000000000000000010); $display(";A 3861");		//(= P1_P3_t    (bv-sdiv P1_P3_r  0b00000000000000000000000000000010))) ;3861
                                                                if ((P1_P3_B == 1'b1)) begin
                                                                    $display(";A 3862");		//(= (bv-comp P1_P3_B  0b1)   0b1)) ;3862
                                                                    P1_P3_t = (P1_P3_t % 32'b00100000000000000000000000000000); $display(";A 3864");		//(= P1_P3_t    (bv-smod P1_P3_t  0b00100000000000000000000000000000))) ;3864
                                                                end
                                                                else begin
                                                                    $display(";A 3863");		//(= (bv-comp P1_P3_B  0b1)   0b0)) ;3863
                                                                end
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 3865");		//(= P1_P3_mf    0b10)) ;3865
                                                                P1_P3_t = ((P1_P3_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 3866");		//(= P1_P3_t    (bv-mul (bv-smod P1_P3_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;3866
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 3867");		//(= P1_P3_mf    0b11)) ;3867
                                                                P1_P3_t = ((P1_P3_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 3868");		//(= P1_P3_t    (bv-mul (bv-smod P1_P3_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;3868
                                                                if ((P1_P3_t > 32'b11111111111111111111111111111111)) begin
                                                                    $display(";A 3869");		//(= (bool-to-bv (bv-gt P1_P3_t  0b11111111111111111111111111111111))   0b1)) ;3869
                                                                    P1_P3_B = 1'b1; $display(";A 3871");		//(= P1_P3_B    0b1)) ;3871
                                                                end
                                                                else begin
                                                                    $display(";A 3870");		//(= (bool-to-bv (bv-gt P1_P3_t  0b11111111111111111111111111111111))   0b0)) ;3870
                                                                    P1_P3_B = 1'b0; $display(";A 3872");		//(= P1_P3_B    0b0)) ;3872
                                                                end
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3873");		//(= (and (/= P1_P3_mf  0b00) (/= P1_P3_mf  0b01) (/= P1_P3_mf  0b10) (/= P1_P3_mf  0b11))   true)) ;3873
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                    case (P1_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 3874");		//(= P1_P3_d    0b00000000000000000000000000000000)) ;3874
                                                                P1_P3_reg0 = P1_P3_t; $display(";A 3875");		//(= P1_P3_reg0    P1_P3_t )) ;3875
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 3876");		//(= P1_P3_d    0b00000000000000000000000000000001)) ;3876
                                                                P1_P3_reg1 = P1_P3_t; $display(";A 3877");		//(= P1_P3_reg1    P1_P3_t )) ;3877
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 3878");		//(= P1_P3_d    0b00000000000000000000000000000010)) ;3878
                                                                P1_P3_reg2 = P1_P3_t; $display(";A 3879");		//(= P1_P3_reg2    P1_P3_t )) ;3879
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 3880");		//(= P1_P3_d    0b00000000000000000000000000000011)) ;3880
                                                                P1_P3_reg3 = P1_P3_t; $display(";A 3881");		//(= P1_P3_reg3    P1_P3_t )) ;3881
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 3882");		//(= (and (/= P1_P3_d  0b00000000000000000000000000000000) (/= P1_P3_d  0b00000000000000000000000000000001) (/= P1_P3_d  0b00000000000000000000000000000010) (/= P1_P3_d  0b00000000000000000000000000000011))   true)) ;3882
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1101 :
                                                begin
                                                    $display(";A 3883");		//(= P1_P3_ff    0b1101)) ;3883
                                                    begin
                                                    end
                                                end
                                            4'b1110 :
                                                begin
                                                    $display(";A 3884");		//(= P1_P3_ff    0b1110)) ;3884
                                                    begin
                                                    end
                                                end
                                            4'b1111 :
                                                begin
                                                    $display(";A 3885");		//(= P1_P3_ff    0b1111)) ;3885
                                                    begin
                                                    end
                                                end
                                        endcase
                                    end
                                    else begin
                                        $display(";A 3552");		//(= (bv-not (bv-comp P1_P3_df  0b00000000000000000000000000000111))   0b0)) ;3552
                                        if ((P1_P3_df == 32'b00000000000000000000000000000111)) begin
                                            $display(";A 3886");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000111)   0b1)) ;3886
                                            case (P1_P3_mf)
                                                2'b00 :
                                                    begin
                                                        $display(";A 3888");		//(= P1_P3_mf    0b00)) ;3888
                                                        P1_P3_m = P1_P3_tail; $display(";A 3889");		//(= P1_P3_m    P1_P3_tail )) ;3889
                                                    end
                                                2'b01 :
                                                    begin
                                                        $display(";A 3890");		//(= P1_P3_mf    0b01)) ;3890
                                                        P1_P3_m = P1_P3_tail; $display(";A 3891");		//(= P1_P3_m    P1_P3_tail )) ;3891
                                                    end
                                                2'b10 :
                                                    begin
                                                        $display(";A 3892");		//(= P1_P3_mf    0b10)) ;3892
                                                        P1_P3_m = ((P1_P3_reg1 % 32'b00000000000100000000000000000000) + (P1_P3_tail % 32'b00000000000100000000000000000000)); $display(";A 3893");		//(= P1_P3_m    (bv-add (bv-smod P1_P3_reg1  0b00000000000100000000000000000000) (bv-smod P1_P3_tail  0b00000000000100000000000000000000)))) ;3893
                                                    end
                                                2'b11 :
                                                    begin
                                                        $display(";A 3894");		//(= P1_P3_mf    0b11)) ;3894
                                                        P1_P3_m = ((P1_P3_reg2 % 32'b00000000000100000000000000000000) + (P1_P3_tail % 32'b00000000000100000000000000000000)); $display(";A 3895");		//(= P1_P3_m    (bv-add (bv-smod P1_P3_reg2  0b00000000000100000000000000000000) (bv-smod P1_P3_tail  0b00000000000100000000000000000000)))) ;3895
                                                    end
                                            endcase
                                            P1_P3_addr <= #1 ((P1_P3_m % 32'sb00000000000000000000000000000010) * 32'sb00000000000000000000000000010100); $display(";A 3896");		//(= P1_P3_addr    (bv-mul (bv-smod P1_P3_m  0b00000000000000000000000000000010) 0b00000000000000000000000000010100))) ;3896
                                            P1_P3_wr <= #1 1'b1; $display(";A 3897");		//(= P1_P3_wr    0b1)) ;3897
                                            P1_P3_datao <= #1 P1_P3_r; $display(";A 3898");		//(= P1_P3_datao    P1_P3_r )) ;3898
                                        end
                                        else begin
                                            $display(";A 3887");		//(= (bv-comp P1_P3_df  0b00000000000000000000000000000111)   0b0)) ;3887
                                        end
                                    end
                                end
                        endcase
                        P1_P3_state = 1'sb0; $display(";A 3899");		//(= P1_P3_state    0b0)) ;3899
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:5810
    always @(posedge P1_P4_reset or posedge P1_P4_clock) begin
        if ((P1_P4_reset == 1'b1)) begin
            P1_P4_MAR = 20'sb00000000000000000000; $display(";A 3902");		//(= P1_P4_MAR    0b00000000000000000000)) ;3902
            P1_P4_MBR = 32'sb00000000000000000000000000000000; $display(";A 3903");		//(= P1_P4_MBR    0b00000000000000000000000000000000)) ;3903
            P1_P4_IR = 32'sb00000000000000000000000000000000; $display(";A 3904");		//(= P1_P4_IR    0b00000000000000000000000000000000)) ;3904
            P1_P4_d = 32'sb00000000000000000000000000000000; $display(";A 3905");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;3905
            P1_P4_r = 32'sb00000000000000000000000000000000; $display(";A 3906");		//(= P1_P4_r    0b00000000000000000000000000000000)) ;3906
            P1_P4_m = 32'sb00000000000000000000000000000000; $display(";A 3907");		//(= P1_P4_m    0b00000000000000000000000000000000)) ;3907
            P1_P4_s = 2'sb00; $display(";A 3908");		//(= P1_P4_s    0b00)) ;3908
            P1_P4_temp = 32'sb00000000000000000000000000000000; $display(";A 3909");		//(= P1_P4_temp    0b00000000000000000000000000000000)) ;3909
            P1_P4_mf = 2'sb00; $display(";A 3910");		//(= P1_P4_mf    0b00)) ;3910
            P1_P4_df = 3'sb000; $display(";A 3911");		//(= P1_P4_df    0b000)) ;3911
            P1_P4_ff = 4'sb0000; $display(";A 3912");		//(= P1_P4_ff    0b0000)) ;3912
            P1_P4_cf = 1'sb0; $display(";A 3913");		//(= P1_P4_cf    0b0)) ;3913
            P1_P4_tail = 20'sb00000000000000000000; $display(";A 3914");		//(= P1_P4_tail    0b00000000000000000000)) ;3914
            P1_P4_B = 1'b0; $display(";A 3915");		//(= P1_P4_B    0b0)) ;3915
            P1_P4_reg0 = 32'sb00000000000000000000000000000000; $display(";A 3916");		//(= P1_P4_reg0    0b00000000000000000000000000000000)) ;3916
            P1_P4_reg1 = 32'sb00000000000000000000000000000000; $display(";A 3917");		//(= P1_P4_reg1    0b00000000000000000000000000000000)) ;3917
            P1_P4_reg2 = 32'sb00000000000000000000000000000000; $display(";A 3918");		//(= P1_P4_reg2    0b00000000000000000000000000000000)) ;3918
            P1_P4_reg3 = 32'sb00000000000000000000000000000000; $display(";A 3919");		//(= P1_P4_reg3    0b00000000000000000000000000000000)) ;3919
            P1_P4_addr <= #1 20'sb00000000000000000000; $display(";A 3920");		//(= P1_P4_addr    0b00000000000000000000)) ;3920
            P1_P4_rd <= #1 1'b0; $display(";A 3921");		//(= P1_P4_rd    0b0)) ;3921
            P1_P4_wr <= #1 1'b0; $display(";A 3922");		//(= P1_P4_wr    0b0)) ;3922
            P1_P4_datao <= #1 32'sb00000000000000000000000000000000; $display(";A 3923");		//(= P1_P4_datao    0b00000000000000000000000000000000)) ;3923
            P1_P4_state = 1'sb0; $display(";A 3924");		//(= P1_P4_state    0b0)) ;3924
        end
        else begin
            P1_P4_rd <= #1 1'b0; $display(";A 3925");		//(= P1_P4_rd    0b0)) ;3925
            P1_P4_wr <= #1 1'b0; $display(";A 3926");		//(= P1_P4_wr    0b0)) ;3926
            case (P1_P4_state)
                1'b0 :
                    begin
                        $display(";A 3927");		//(= P1_P4_state    0b0)) ;3927
                        P1_P4_MAR = (P1_P4_reg3 % 32'b00000000000100000000000000000000); $display(";A 3928");		//(= P1_P4_MAR    (bv-smod P1_P4_reg3  0b00000000000100000000000000000000))) ;3928
                        P1_P4_addr <= #1 P1_P4_MAR; $display(";A 3929");		//(= P1_P4_addr    P1_P4_MAR )) ;3929
                        P1_P4_rd <= #1 1'b1; $display(";A 3930");		//(= P1_P4_rd    0b1)) ;3930
                        P1_P4_MBR = P1_P4_datai; $display(";A 3931");		//(= P1_P4_MBR    P1_P4_datai )) ;3931
                        P1_P4_IR = P1_P4_MBR; $display(";A 3932");		//(= P1_P4_IR    P1_P4_MBR )) ;3932
                        P1_P4_state = 1'sb1; $display(";A 3933");		//(= P1_P4_state    0b1)) ;3933
                    end
                1'b1 :
                    begin
                        $display(";A 3934");		//(= P1_P4_state    0b1)) ;3934
                        if ((P1_P4_IR < 32'sb00000000000000000000000000000000)) begin
                            $display(";A 3935");		//(= (bool-to-bv (bv-slt P1_P4_IR  0b00000000000000000000000000000000))   0b1)) ;3935
                            P1_P4_IR = (-P1_P4_IR); $display(";A 3937");		//(= P1_P4_IR    (bv-neg P1_P4_IR ))) ;3937
                        end
                        else begin
                            $display(";A 3936");		//(= (bool-to-bv (bv-slt P1_P4_IR  0b00000000000000000000000000000000))   0b0)) ;3936
                        end
                        P1_P4_mf = ((P1_P4_IR / 32'b00001000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 3938");		//(= P1_P4_mf    (bv-smod (bv-sdiv P1_P4_IR  0b00001000000000000000000000000000) 0b00000000000000000000000000000100))) ;3938
                        P1_P4_df = ((P1_P4_IR / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000000001000); $display(";A 3939");		//(= P1_P4_df    (bv-smod (bv-sdiv P1_P4_IR  0b00000001000000000000000000000000) 0b00000000000000000000000000001000))) ;3939
                        P1_P4_ff = ((P1_P4_IR / 32'b00000000000010000000000000000000) % 32'b00000000000000000000000000010000); $display(";A 3940");		//(= P1_P4_ff    (bv-smod (bv-sdiv P1_P4_IR  0b00000000000010000000000000000000) 0b00000000000000000000000000010000))) ;3940
                        P1_P4_cf = ((P1_P4_IR / 32'b00000000100000000000000000000000) % 32'b00000000000000000000000000000010); $display(";A 3941");		//(= P1_P4_cf    (bv-smod (bv-sdiv P1_P4_IR  0b00000000100000000000000000000000) 0b00000000000000000000000000000010))) ;3941
                        P1_P4_tail = (P1_P4_IR % 32'b00000000000100000000000000000000); $display(";A 3942");		//(= P1_P4_tail    (bv-smod P1_P4_IR  0b00000000000100000000000000000000))) ;3942
                        P1_P4_reg3 = ((P1_P4_reg3 % 32'b00100000000000000000000000000000) + 32'b00000000000000000000000000001000); $display(";A 3943");		//(= P1_P4_reg3    (bv-add (bv-smod P1_P4_reg3  0b00100000000000000000000000000000) 0b00000000000000000000000000001000))) ;3943
                        P1_P4_s = ((P1_P4_IR / 32'b00100000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 3944");		//(= P1_P4_s    (bv-smod (bv-sdiv P1_P4_IR  0b00100000000000000000000000000000) 0b00000000000000000000000000000100))) ;3944
                        case (P1_P4_s)
                            2'b00 :
                                begin
                                    $display(";A 3945");		//(= P1_P4_s    0b00)) ;3945
                                    P1_P4_r = P1_P4_reg0; $display(";A 3946");		//(= P1_P4_r    P1_P4_reg0 )) ;3946
                                end
                            2'b01 :
                                begin
                                    $display(";A 3947");		//(= P1_P4_s    0b01)) ;3947
                                    P1_P4_r = P1_P4_reg1; $display(";A 3948");		//(= P1_P4_r    P1_P4_reg1 )) ;3948
                                end
                            2'b10 :
                                begin
                                    $display(";A 3949");		//(= P1_P4_s    0b10)) ;3949
                                    P1_P4_r = P1_P4_reg2; $display(";A 3950");		//(= P1_P4_r    P1_P4_reg2 )) ;3950
                                end
                            2'b11 :
                                begin
                                    $display(";A 3951");		//(= P1_P4_s    0b11)) ;3951
                                    P1_P4_r = P1_P4_reg3; $display(";A 3952");		//(= P1_P4_r    P1_P4_reg3 )) ;3952
                                end
                        endcase
                        case (P1_P4_cf)
                            1'b1 :
                                begin
                                    $display(";A 3953");		//(= P1_P4_cf    0b1)) ;3953
                                    case (P1_P4_mf)
                                        2'b00 :
                                            begin
                                                $display(";A 3954");		//(= P1_P4_mf    0b00)) ;3954
                                                P1_P4_m = P1_P4_tail; $display(";A 3955");		//(= P1_P4_m    P1_P4_tail )) ;3955
                                            end
                                        2'b01 :
                                            begin
                                                $display(";A 3956");		//(= P1_P4_mf    0b01)) ;3956
                                                P1_P4_m = P1_P4_datai; $display(";A 3957");		//(= P1_P4_m    P1_P4_datai )) ;3957
                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 3958");		//(= P1_P4_addr    P1_P4_tail )) ;3958
                                                P1_P4_rd <= #1 1'b1; $display(";A 3959");		//(= P1_P4_rd    0b1)) ;3959
                                            end
                                        2'b10 :
                                            begin
                                                $display(";A 3960");		//(= P1_P4_mf    0b10)) ;3960
                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 3961");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;3961
                                                P1_P4_rd <= #1 1'b1; $display(";A 3962");		//(= P1_P4_rd    0b1)) ;3962
                                                P1_P4_m = P1_P4_datai; $display(";A 3963");		//(= P1_P4_m    P1_P4_datai )) ;3963
                                            end
                                        2'b11 :
                                            begin
                                                $display(";A 3964");		//(= P1_P4_mf    0b11)) ;3964
                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 3965");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;3965
                                                P1_P4_rd <= #1 1'b1; $display(";A 3966");		//(= P1_P4_rd    0b1)) ;3966
                                                P1_P4_m = P1_P4_datai; $display(";A 3967");		//(= P1_P4_m    P1_P4_datai )) ;3967
                                            end
                                    endcase
                                    case (P1_P4_ff)
                                        4'b0000 :
                                            begin
                                                $display(";A 3968");		//(= P1_P4_ff    0b0000)) ;3968
                                                if ((P1_P4_r < P1_P4_m)) begin
                                                    $display(";A 3969");		//(= (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))   0b1)) ;3969
                                                    P1_P4_B = 1'b1; $display(";A 3971");		//(= P1_P4_B    0b1)) ;3971
                                                end
                                                else begin
                                                    $display(";A 3970");		//(= (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))   0b0)) ;3970
                                                    P1_P4_B = 1'b0; $display(";A 3972");		//(= P1_P4_B    0b0)) ;3972
                                                end
                                            end
                                        4'b0001 :
                                            begin
                                                $display(";A 3973");		//(= P1_P4_ff    0b0001)) ;3973
                                                if ((~(P1_P4_r < P1_P4_m))) begin
                                                    $display(";A 3974");		//(= (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )))   0b1)) ;3974
                                                    P1_P4_B = 1'b1; $display(";A 3976");		//(= P1_P4_B    0b1)) ;3976
                                                end
                                                else begin
                                                    $display(";A 3975");		//(= (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )))   0b0)) ;3975
                                                    P1_P4_B = 1'b0; $display(";A 3977");		//(= P1_P4_B    0b0)) ;3977
                                                end
                                            end
                                        4'b0010 :
                                            begin
                                                $display(";A 3978");		//(= P1_P4_ff    0b0010)) ;3978
                                                if ((P1_P4_r == P1_P4_m)) begin
                                                    $display(";A 3979");		//(= (bv-comp P1_P4_r  P1_P4_m )   0b1)) ;3979
                                                    P1_P4_B = 1'b1; $display(";A 3981");		//(= P1_P4_B    0b1)) ;3981
                                                end
                                                else begin
                                                    $display(";A 3980");		//(= (bv-comp P1_P4_r  P1_P4_m )   0b0)) ;3980
                                                    P1_P4_B = 1'b0; $display(";A 3982");		//(= P1_P4_B    0b0)) ;3982
                                                end
                                            end
                                        4'b0011 :
                                            begin
                                                $display(";A 3983");		//(= P1_P4_ff    0b0011)) ;3983
                                                if ((~(P1_P4_r == P1_P4_m))) begin
                                                    $display(";A 3984");		//(= (bv-not (bv-comp P1_P4_r  P1_P4_m ))   0b1)) ;3984
                                                    P1_P4_B = 1'b1; $display(";A 3986");		//(= P1_P4_B    0b1)) ;3986
                                                end
                                                else begin
                                                    $display(";A 3985");		//(= (bv-not (bv-comp P1_P4_r  P1_P4_m ))   0b0)) ;3985
                                                    P1_P4_B = 1'b0; $display(";A 3987");		//(= P1_P4_B    0b0)) ;3987
                                                end
                                            end
                                        4'b0100 :
                                            begin
                                                $display(";A 3988");		//(= P1_P4_ff    0b0100)) ;3988
                                                if ((~(P1_P4_r > P1_P4_m))) begin
                                                    $display(";A 3989");		//(= (bv-not (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m )))   0b1)) ;3989
                                                    P1_P4_B = 1'b1; $display(";A 3991");		//(= P1_P4_B    0b1)) ;3991
                                                end
                                                else begin
                                                    $display(";A 3990");		//(= (bv-not (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m )))   0b0)) ;3990
                                                    P1_P4_B = 1'b0; $display(";A 3992");		//(= P1_P4_B    0b0)) ;3992
                                                end
                                            end
                                        4'b0101 :
                                            begin
                                                $display(";A 3993");		//(= P1_P4_ff    0b0101)) ;3993
                                                if ((P1_P4_r > P1_P4_m)) begin
                                                    $display(";A 3994");		//(= (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m ))   0b1)) ;3994
                                                    P1_P4_B = 1'b1; $display(";A 3996");		//(= P1_P4_B    0b1)) ;3996
                                                end
                                                else begin
                                                    $display(";A 3995");		//(= (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m ))   0b0)) ;3995
                                                    P1_P4_B = 1'b0; $display(";A 3997");		//(= P1_P4_B    0b0)) ;3997
                                                end
                                            end
                                        4'b0110 :
                                            begin
                                                $display(";A 3998");		//(= P1_P4_ff    0b0110)) ;3998
                                                if ((P1_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 3999");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b1)) ;3999
                                                    P1_P4_r = (P1_P4_r - 32'b00000000000000000000000000000000); $display(";A 4001");		//(= P1_P4_r    (bv-sub P1_P4_r  0b00000000000000000000000000000000))) ;4001
                                                end
                                                else begin
                                                    $display(";A 4000");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b0)) ;4000
                                                end
                                                if ((P1_P4_r < P1_P4_m)) begin
                                                    $display(";A 4002");		//(= (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))   0b1)) ;4002
                                                    P1_P4_B = 1'b1; $display(";A 4004");		//(= P1_P4_B    0b1)) ;4004
                                                end
                                                else begin
                                                    $display(";A 4003");		//(= (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))   0b0)) ;4003
                                                    P1_P4_B = 1'b0; $display(";A 4005");		//(= P1_P4_B    0b0)) ;4005
                                                end
                                            end
                                        4'b0111 :
                                            begin
                                                $display(";A 4006");		//(= P1_P4_ff    0b0111)) ;4006
                                                if ((P1_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 4007");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b1)) ;4007
                                                    P1_P4_r = (P1_P4_r - 32'b00000000000000000000000000000000); $display(";A 4009");		//(= P1_P4_r    (bv-sub P1_P4_r  0b00000000000000000000000000000000))) ;4009
                                                end
                                                else begin
                                                    $display(";A 4008");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b0)) ;4008
                                                end
                                                if ((~(P1_P4_r < P1_P4_m))) begin
                                                    $display(";A 4010");		//(= (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )))   0b1)) ;4010
                                                    P1_P4_B = 1'b1; $display(";A 4012");		//(= P1_P4_B    0b1)) ;4012
                                                end
                                                else begin
                                                    $display(";A 4011");		//(= (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )))   0b0)) ;4011
                                                    P1_P4_B = 1'b0; $display(";A 4013");		//(= P1_P4_B    0b0)) ;4013
                                                end
                                            end
                                        4'b1000 :
                                            begin
                                                $display(";A 4014");		//(= P1_P4_ff    0b1000)) ;4014
                                                if (((P1_P4_r < P1_P4_m) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4015");		//(= (bv-or (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b1)) ;4015
                                                    P1_P4_B = 1'b1; $display(";A 4017");		//(= P1_P4_B    0b1)) ;4017
                                                end
                                                else begin
                                                    $display(";A 4016");		//(= (bv-or (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b0)) ;4016
                                                    P1_P4_B = 1'b0; $display(";A 4018");		//(= P1_P4_B    0b0)) ;4018
                                                end
                                            end
                                        4'b1001 :
                                            begin
                                                $display(";A 4019");		//(= P1_P4_ff    0b1001)) ;4019
                                                if (((~(P1_P4_r < P1_P4_m)) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4020");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))) (bv-comp P1_P4_B  0b1))   0b1)) ;4020
                                                    P1_P4_B = 1'b1; $display(";A 4022");		//(= P1_P4_B    0b1)) ;4022
                                                end
                                                else begin
                                                    $display(";A 4021");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))) (bv-comp P1_P4_B  0b1))   0b0)) ;4021
                                                    P1_P4_B = 1'b0; $display(";A 4023");		//(= P1_P4_B    0b0)) ;4023
                                                end
                                            end
                                        4'b1010 :
                                            begin
                                                $display(";A 4024");		//(= P1_P4_ff    0b1010)) ;4024
                                                if (((P1_P4_r == P1_P4_m) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4025");		//(= (bv-or (bv-comp P1_P4_r  P1_P4_m ) (bv-comp P1_P4_B  0b1))   0b1)) ;4025
                                                    P1_P4_B = 1'b1; $display(";A 4027");		//(= P1_P4_B    0b1)) ;4027
                                                end
                                                else begin
                                                    $display(";A 4026");		//(= (bv-or (bv-comp P1_P4_r  P1_P4_m ) (bv-comp P1_P4_B  0b1))   0b0)) ;4026
                                                    P1_P4_B = 1'b0; $display(";A 4028");		//(= P1_P4_B    0b0)) ;4028
                                                end
                                            end
                                        4'b1011 :
                                            begin
                                                $display(";A 4029");		//(= P1_P4_ff    0b1011)) ;4029
                                                if (((~(P1_P4_r == P1_P4_m)) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4030");		//(= (bv-or (bv-not (bv-comp P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b1)) ;4030
                                                    P1_P4_B = 1'b1; $display(";A 4032");		//(= P1_P4_B    0b1)) ;4032
                                                end
                                                else begin
                                                    $display(";A 4031");		//(= (bv-or (bv-not (bv-comp P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b0)) ;4031
                                                    P1_P4_B = 1'b0; $display(";A 4033");		//(= P1_P4_B    0b0)) ;4033
                                                end
                                            end
                                        4'b1100 :
                                            begin
                                                $display(";A 4034");		//(= P1_P4_ff    0b1100)) ;4034
                                                if (((~(P1_P4_r > P1_P4_m)) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4035");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m ))) (bv-comp P1_P4_B  0b1))   0b1)) ;4035
                                                    P1_P4_B = 1'b1; $display(";A 4037");		//(= P1_P4_B    0b1)) ;4037
                                                end
                                                else begin
                                                    $display(";A 4036");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m ))) (bv-comp P1_P4_B  0b1))   0b0)) ;4036
                                                    P1_P4_B = 1'b0; $display(";A 4038");		//(= P1_P4_B    0b0)) ;4038
                                                end
                                            end
                                        4'b1101 :
                                            begin
                                                $display(";A 4039");		//(= P1_P4_ff    0b1101)) ;4039
                                                if (((P1_P4_r > P1_P4_m) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4040");		//(= (bv-or (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b1)) ;4040
                                                    P1_P4_B = 1'b1; $display(";A 4042");		//(= P1_P4_B    0b1)) ;4042
                                                end
                                                else begin
                                                    $display(";A 4041");		//(= (bv-or (bool-to-bv (bv-sgt P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b0)) ;4041
                                                    P1_P4_B = 1'b0; $display(";A 4043");		//(= P1_P4_B    0b0)) ;4043
                                                end
                                            end
                                        4'b1110 :
                                            begin
                                                $display(";A 4044");		//(= P1_P4_ff    0b1110)) ;4044
                                                if ((P1_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 4045");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b1)) ;4045
                                                    P1_P4_r = (P1_P4_r - 32'b00000000000000000000000000000000); $display(";A 4047");		//(= P1_P4_r    (bv-sub P1_P4_r  0b00000000000000000000000000000000))) ;4047
                                                end
                                                else begin
                                                    $display(";A 4046");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b0)) ;4046
                                                end
                                                if (((P1_P4_r < P1_P4_m) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4048");		//(= (bv-or (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b1)) ;4048
                                                    P1_P4_B = 1'b1; $display(";A 4050");		//(= P1_P4_B    0b1)) ;4050
                                                end
                                                else begin
                                                    $display(";A 4049");		//(= (bv-or (bool-to-bv (bv-slt P1_P4_r  P1_P4_m )) (bv-comp P1_P4_B  0b1))   0b0)) ;4049
                                                    P1_P4_B = 1'b0; $display(";A 4051");		//(= P1_P4_B    0b0)) ;4051
                                                end
                                            end
                                        4'b1111 :
                                            begin
                                                $display(";A 4052");		//(= P1_P4_ff    0b1111)) ;4052
                                                if ((P1_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 4053");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b1)) ;4053
                                                    P1_P4_r = (P1_P4_r - 32'b00000000000000000000000000000000); $display(";A 4055");		//(= P1_P4_r    (bv-sub P1_P4_r  0b00000000000000000000000000000000))) ;4055
                                                end
                                                else begin
                                                    $display(";A 4054");		//(= (bool-to-bv (bv-gt P1_P4_r  0b11111111111111111111111111111111))   0b0)) ;4054
                                                end
                                                if (((~(P1_P4_r < P1_P4_m)) | (P1_P4_B == 1'b1))) begin
                                                    $display(";A 4056");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))) (bv-comp P1_P4_B  0b1))   0b1)) ;4056
                                                    P1_P4_B = 1'b1; $display(";A 4058");		//(= P1_P4_B    0b1)) ;4058
                                                end
                                                else begin
                                                    $display(";A 4057");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P1_P4_r  P1_P4_m ))) (bv-comp P1_P4_B  0b1))   0b0)) ;4057
                                                    P1_P4_B = 1'b0; $display(";A 4059");		//(= P1_P4_B    0b0)) ;4059
                                                end
                                            end
                                    endcase
                                end
                            1'b0 :
                                begin
                                    $display(";A 4060");		//(= P1_P4_cf    0b0)) ;4060
                                    if ((~(P1_P4_df == 32'b00000000000000000000000000000111))) begin
                                        $display(";A 4061");		//(= (bv-not (bv-comp P1_P4_df  0b00000000000000000000000000000111))   0b1)) ;4061
                                        if ((P1_P4_df == 32'b00000000000000000000000000000101)) begin
                                            $display(";A 4063");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000101)   0b1)) ;4063
                                            if (((~P1_P4_B) == 1'b1)) begin
                                                $display(";A 4065");		//(= (bv-comp (bv-not P1_P4_B ) 0b1)   0b1)) ;4065
                                                P1_P4_d = 32'sb00000000000000000000000000000011; $display(";A 4067");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4067
                                            end
                                            else begin
                                                $display(";A 4066");		//(= (bv-comp (bv-not P1_P4_B ) 0b1)   0b0)) ;4066
                                            end
                                        end
                                        else begin
                                            $display(";A 4064");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000101)   0b0)) ;4064
                                            if ((P1_P4_df == 32'b00000000000000000000000000000100)) begin
                                                $display(";A 4068");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000100)   0b1)) ;4068
                                                if ((P1_P4_B == 1'b1)) begin
                                                    $display(";A 4070");		//(= (bv-comp P1_P4_B  0b1)   0b1)) ;4070
                                                    P1_P4_d = 32'sb00000000000000000000000000000011; $display(";A 4072");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4072
                                                end
                                                else begin
                                                    $display(";A 4071");		//(= (bv-comp P1_P4_B  0b1)   0b0)) ;4071
                                                end
                                            end
                                            else begin
                                                $display(";A 4069");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000100)   0b0)) ;4069
                                                if ((P1_P4_df == 32'b00000000000000000000000000000011)) begin
                                                    $display(";A 4073");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000011)   0b1)) ;4073
                                                    P1_P4_d = 32'sb00000000000000000000000000000011; $display(";A 4075");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4075
                                                end
                                                else begin
                                                    $display(";A 4074");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000011)   0b0)) ;4074
                                                    if ((P1_P4_df == 32'b00000000000000000000000000000010)) begin
                                                        $display(";A 4076");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000010)   0b1)) ;4076
                                                        P1_P4_d = 32'sb00000000000000000000000000000010; $display(";A 4078");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4078
                                                    end
                                                    else begin
                                                        $display(";A 4077");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000010)   0b0)) ;4077
                                                        if ((P1_P4_df == 32'b00000000000000000000000000000001)) begin
                                                            $display(";A 4079");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000001)   0b1)) ;4079
                                                            P1_P4_d = 32'sb00000000000000000000000000000001; $display(";A 4081");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4081
                                                        end
                                                        else begin
                                                            $display(";A 4080");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000001)   0b0)) ;4080
                                                            if ((P1_P4_df == 32'b00000000000000000000000000000000)) begin
                                                                $display(";A 4082");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000000)   0b1)) ;4082
                                                                P1_P4_d = 32'sb00000000000000000000000000000000; $display(";A 4084");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4084
                                                            end
                                                            else begin
                                                                $display(";A 4083");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000000)   0b0)) ;4083
                                                            end
                                                        end
                                                    end
                                                end
                                            end
                                        end
                                        case (P1_P4_ff)
                                            4'b0000 :
                                                begin
                                                    $display(";A 4085");		//(= P1_P4_ff    0b0000)) ;4085
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4086");		//(= P1_P4_mf    0b00)) ;4086
                                                                P1_P4_m = P1_P4_tail; $display(";A 4087");		//(= P1_P4_m    P1_P4_tail )) ;4087
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4088");		//(= P1_P4_mf    0b01)) ;4088
                                                                P1_P4_m = P1_P4_datai; $display(";A 4089");		//(= P1_P4_m    P1_P4_datai )) ;4089
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4090");		//(= P1_P4_addr    P1_P4_tail )) ;4090
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4091");		//(= P1_P4_rd    0b1)) ;4091
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4092");		//(= P1_P4_mf    0b10)) ;4092
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4093");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4093
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4094");		//(= P1_P4_rd    0b1)) ;4094
                                                                P1_P4_m = P1_P4_datai; $display(";A 4095");		//(= P1_P4_m    P1_P4_datai )) ;4095
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4096");		//(= P1_P4_mf    0b11)) ;4096
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4097");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4097
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4098");		//(= P1_P4_rd    0b1)) ;4098
                                                                P1_P4_m = P1_P4_datai; $display(";A 4099");		//(= P1_P4_m    P1_P4_datai )) ;4099
                                                            end
                                                    endcase
                                                    P1_P4_t = 32'sb00000000000000000000000000000000; $display(";A 4100");		//(= P1_P4_t    0b00000000000000000000000000000000)) ;4100
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4101");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4101
                                                                P1_P4_reg0 = (P1_P4_t - P1_P4_m); $display(";A 4102");		//(= P1_P4_reg0    (bv-sub P1_P4_t  P1_P4_m ))) ;4102
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4103");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4103
                                                                P1_P4_reg1 = (P1_P4_t - P1_P4_m); $display(";A 4104");		//(= P1_P4_reg1    (bv-sub P1_P4_t  P1_P4_m ))) ;4104
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4105");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4105
                                                                P1_P4_reg2 = (P1_P4_t - P1_P4_m); $display(";A 4106");		//(= P1_P4_reg2    (bv-sub P1_P4_t  P1_P4_m ))) ;4106
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4107");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4107
                                                                P1_P4_reg3 = (P1_P4_t - P1_P4_m); $display(";A 4108");		//(= P1_P4_reg3    (bv-sub P1_P4_t  P1_P4_m ))) ;4108
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4109");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4109
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0001 :
                                                begin
                                                    $display(";A 4110");		//(= P1_P4_ff    0b0001)) ;4110
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4111");		//(= P1_P4_mf    0b00)) ;4111
                                                                P1_P4_m = P1_P4_tail; $display(";A 4112");		//(= P1_P4_m    P1_P4_tail )) ;4112
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4113");		//(= P1_P4_mf    0b01)) ;4113
                                                                P1_P4_m = P1_P4_datai; $display(";A 4114");		//(= P1_P4_m    P1_P4_datai )) ;4114
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4115");		//(= P1_P4_addr    P1_P4_tail )) ;4115
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4116");		//(= P1_P4_rd    0b1)) ;4116
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4117");		//(= P1_P4_mf    0b10)) ;4117
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4118");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4118
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4119");		//(= P1_P4_rd    0b1)) ;4119
                                                                P1_P4_m = P1_P4_datai; $display(";A 4120");		//(= P1_P4_m    P1_P4_datai )) ;4120
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4121");		//(= P1_P4_mf    0b11)) ;4121
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4122");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4122
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4123");		//(= P1_P4_rd    0b1)) ;4123
                                                                P1_P4_m = P1_P4_datai; $display(";A 4124");		//(= P1_P4_m    P1_P4_datai )) ;4124
                                                            end
                                                    endcase
                                                    P1_P4_reg2 = P1_P4_reg3; $display(";A 4125");		//(= P1_P4_reg2    P1_P4_reg3 )) ;4125
                                                    P1_P4_reg3 = P1_P4_m; $display(";A 4126");		//(= P1_P4_reg3    P1_P4_m )) ;4126
                                                end
                                            4'b0010 :
                                                begin
                                                    $display(";A 4127");		//(= P1_P4_ff    0b0010)) ;4127
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4128");		//(= P1_P4_mf    0b00)) ;4128
                                                                P1_P4_m = P1_P4_tail; $display(";A 4129");		//(= P1_P4_m    P1_P4_tail )) ;4129
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4130");		//(= P1_P4_mf    0b01)) ;4130
                                                                P1_P4_m = P1_P4_datai; $display(";A 4131");		//(= P1_P4_m    P1_P4_datai )) ;4131
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4132");		//(= P1_P4_addr    P1_P4_tail )) ;4132
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4133");		//(= P1_P4_rd    0b1)) ;4133
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4134");		//(= P1_P4_mf    0b10)) ;4134
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4135");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4135
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4136");		//(= P1_P4_rd    0b1)) ;4136
                                                                P1_P4_m = P1_P4_datai; $display(";A 4137");		//(= P1_P4_m    P1_P4_datai )) ;4137
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4138");		//(= P1_P4_mf    0b11)) ;4138
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4139");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4139
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4140");		//(= P1_P4_rd    0b1)) ;4140
                                                                P1_P4_m = P1_P4_datai; $display(";A 4141");		//(= P1_P4_m    P1_P4_datai )) ;4141
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4142");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4142
                                                                P1_P4_reg0 = P1_P4_m; $display(";A 4143");		//(= P1_P4_reg0    P1_P4_m )) ;4143
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4144");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4144
                                                                P1_P4_reg1 = P1_P4_m; $display(";A 4145");		//(= P1_P4_reg1    P1_P4_m )) ;4145
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4146");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4146
                                                                P1_P4_reg2 = P1_P4_m; $display(";A 4147");		//(= P1_P4_reg2    P1_P4_m )) ;4147
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4148");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4148
                                                                P1_P4_reg3 = P1_P4_m; $display(";A 4149");		//(= P1_P4_reg3    P1_P4_m )) ;4149
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4150");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4150
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0011 :
                                                begin
                                                    $display(";A 4151");		//(= P1_P4_ff    0b0011)) ;4151
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4152");		//(= P1_P4_mf    0b00)) ;4152
                                                                P1_P4_m = P1_P4_tail; $display(";A 4153");		//(= P1_P4_m    P1_P4_tail )) ;4153
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4154");		//(= P1_P4_mf    0b01)) ;4154
                                                                P1_P4_m = P1_P4_datai; $display(";A 4155");		//(= P1_P4_m    P1_P4_datai )) ;4155
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4156");		//(= P1_P4_addr    P1_P4_tail )) ;4156
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4157");		//(= P1_P4_rd    0b1)) ;4157
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4158");		//(= P1_P4_mf    0b10)) ;4158
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4159");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4159
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4160");		//(= P1_P4_rd    0b1)) ;4160
                                                                P1_P4_m = P1_P4_datai; $display(";A 4161");		//(= P1_P4_m    P1_P4_datai )) ;4161
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4162");		//(= P1_P4_mf    0b11)) ;4162
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4163");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4163
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4164");		//(= P1_P4_rd    0b1)) ;4164
                                                                P1_P4_m = P1_P4_datai; $display(";A 4165");		//(= P1_P4_m    P1_P4_datai )) ;4165
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4166");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4166
                                                                P1_P4_reg0 = P1_P4_m; $display(";A 4167");		//(= P1_P4_reg0    P1_P4_m )) ;4167
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4168");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4168
                                                                P1_P4_reg1 = P1_P4_m; $display(";A 4169");		//(= P1_P4_reg1    P1_P4_m )) ;4169
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4170");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4170
                                                                P1_P4_reg2 = P1_P4_m; $display(";A 4171");		//(= P1_P4_reg2    P1_P4_m )) ;4171
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4172");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4172
                                                                P1_P4_reg3 = P1_P4_m; $display(";A 4173");		//(= P1_P4_reg3    P1_P4_m )) ;4173
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4174");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4174
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0100 :
                                                begin
                                                    $display(";A 4175");		//(= P1_P4_ff    0b0100)) ;4175
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4176");		//(= P1_P4_mf    0b00)) ;4176
                                                                P1_P4_m = P1_P4_tail; $display(";A 4177");		//(= P1_P4_m    P1_P4_tail )) ;4177
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4178");		//(= P1_P4_mf    0b01)) ;4178
                                                                P1_P4_m = P1_P4_datai; $display(";A 4179");		//(= P1_P4_m    P1_P4_datai )) ;4179
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4180");		//(= P1_P4_addr    P1_P4_tail )) ;4180
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4181");		//(= P1_P4_rd    0b1)) ;4181
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4182");		//(= P1_P4_mf    0b10)) ;4182
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4183");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4183
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4184");		//(= P1_P4_rd    0b1)) ;4184
                                                                P1_P4_m = P1_P4_datai; $display(";A 4185");		//(= P1_P4_m    P1_P4_datai )) ;4185
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4186");		//(= P1_P4_mf    0b11)) ;4186
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4187");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4187
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4188");		//(= P1_P4_rd    0b1)) ;4188
                                                                P1_P4_m = P1_P4_datai; $display(";A 4189");		//(= P1_P4_m    P1_P4_datai )) ;4189
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4190");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4190
                                                                P1_P4_reg0 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4191");		//(= P1_P4_reg0    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4191
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4192");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4192
                                                                P1_P4_reg1 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4193");		//(= P1_P4_reg1    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4193
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4194");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4194
                                                                P1_P4_reg2 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4195");		//(= P1_P4_reg2    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4195
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4196");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4196
                                                                P1_P4_reg3 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4197");		//(= P1_P4_reg3    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4197
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4198");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4198
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0101 :
                                                begin
                                                    $display(";A 4199");		//(= P1_P4_ff    0b0101)) ;4199
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4200");		//(= P1_P4_mf    0b00)) ;4200
                                                                P1_P4_m = P1_P4_tail; $display(";A 4201");		//(= P1_P4_m    P1_P4_tail )) ;4201
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4202");		//(= P1_P4_mf    0b01)) ;4202
                                                                P1_P4_m = P1_P4_datai; $display(";A 4203");		//(= P1_P4_m    P1_P4_datai )) ;4203
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4204");		//(= P1_P4_addr    P1_P4_tail )) ;4204
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4205");		//(= P1_P4_rd    0b1)) ;4205
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4206");		//(= P1_P4_mf    0b10)) ;4206
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4207");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4207
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4208");		//(= P1_P4_rd    0b1)) ;4208
                                                                P1_P4_m = P1_P4_datai; $display(";A 4209");		//(= P1_P4_m    P1_P4_datai )) ;4209
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4210");		//(= P1_P4_mf    0b11)) ;4210
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4211");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4211
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4212");		//(= P1_P4_rd    0b1)) ;4212
                                                                P1_P4_m = P1_P4_datai; $display(";A 4213");		//(= P1_P4_m    P1_P4_datai )) ;4213
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4214");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4214
                                                                P1_P4_reg0 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4215");		//(= P1_P4_reg0    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4215
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4216");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4216
                                                                P1_P4_reg1 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4217");		//(= P1_P4_reg1    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4217
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4218");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4218
                                                                P1_P4_reg2 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4219");		//(= P1_P4_reg2    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4219
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4220");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4220
                                                                P1_P4_reg3 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4221");		//(= P1_P4_reg3    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4221
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4222");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4222
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0110 :
                                                begin
                                                    $display(";A 4223");		//(= P1_P4_ff    0b0110)) ;4223
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4224");		//(= P1_P4_mf    0b00)) ;4224
                                                                P1_P4_m = P1_P4_tail; $display(";A 4225");		//(= P1_P4_m    P1_P4_tail )) ;4225
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4226");		//(= P1_P4_mf    0b01)) ;4226
                                                                P1_P4_m = P1_P4_datai; $display(";A 4227");		//(= P1_P4_m    P1_P4_datai )) ;4227
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4228");		//(= P1_P4_addr    P1_P4_tail )) ;4228
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4229");		//(= P1_P4_rd    0b1)) ;4229
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4230");		//(= P1_P4_mf    0b10)) ;4230
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4231");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4231
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4232");		//(= P1_P4_rd    0b1)) ;4232
                                                                P1_P4_m = P1_P4_datai; $display(";A 4233");		//(= P1_P4_m    P1_P4_datai )) ;4233
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4234");		//(= P1_P4_mf    0b11)) ;4234
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4235");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4235
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4236");		//(= P1_P4_rd    0b1)) ;4236
                                                                P1_P4_m = P1_P4_datai; $display(";A 4237");		//(= P1_P4_m    P1_P4_datai )) ;4237
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4238");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4238
                                                                P1_P4_reg0 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4239");		//(= P1_P4_reg0    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4239
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4240");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4240
                                                                P1_P4_reg1 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4241");		//(= P1_P4_reg1    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4241
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4242");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4242
                                                                P1_P4_reg2 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4243");		//(= P1_P4_reg2    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4243
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4244");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4244
                                                                P1_P4_reg3 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4245");		//(= P1_P4_reg3    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4245
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4246");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4246
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0111 :
                                                begin
                                                    $display(";A 4247");		//(= P1_P4_ff    0b0111)) ;4247
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4248");		//(= P1_P4_mf    0b00)) ;4248
                                                                P1_P4_m = P1_P4_tail; $display(";A 4249");		//(= P1_P4_m    P1_P4_tail )) ;4249
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4250");		//(= P1_P4_mf    0b01)) ;4250
                                                                P1_P4_m = P1_P4_datai; $display(";A 4251");		//(= P1_P4_m    P1_P4_datai )) ;4251
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4252");		//(= P1_P4_addr    P1_P4_tail )) ;4252
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4253");		//(= P1_P4_rd    0b1)) ;4253
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4254");		//(= P1_P4_mf    0b10)) ;4254
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4255");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4255
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4256");		//(= P1_P4_rd    0b1)) ;4256
                                                                P1_P4_m = P1_P4_datai; $display(";A 4257");		//(= P1_P4_m    P1_P4_datai )) ;4257
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4258");		//(= P1_P4_mf    0b11)) ;4258
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4259");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4259
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4260");		//(= P1_P4_rd    0b1)) ;4260
                                                                P1_P4_m = P1_P4_datai; $display(";A 4261");		//(= P1_P4_m    P1_P4_datai )) ;4261
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4262");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4262
                                                                P1_P4_reg0 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4263");		//(= P1_P4_reg0    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4263
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4264");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4264
                                                                P1_P4_reg1 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4265");		//(= P1_P4_reg1    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4265
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4266");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4266
                                                                P1_P4_reg2 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4267");		//(= P1_P4_reg2    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4267
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4268");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4268
                                                                P1_P4_reg3 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4269");		//(= P1_P4_reg3    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4269
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4270");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4270
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1000 :
                                                begin
                                                    $display(";A 4271");		//(= P1_P4_ff    0b1000)) ;4271
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4272");		//(= P1_P4_mf    0b00)) ;4272
                                                                P1_P4_m = P1_P4_tail; $display(";A 4273");		//(= P1_P4_m    P1_P4_tail )) ;4273
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4274");		//(= P1_P4_mf    0b01)) ;4274
                                                                P1_P4_m = P1_P4_datai; $display(";A 4275");		//(= P1_P4_m    P1_P4_datai )) ;4275
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4276");		//(= P1_P4_addr    P1_P4_tail )) ;4276
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4277");		//(= P1_P4_rd    0b1)) ;4277
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4278");		//(= P1_P4_mf    0b10)) ;4278
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4279");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4279
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4280");		//(= P1_P4_rd    0b1)) ;4280
                                                                P1_P4_m = P1_P4_datai; $display(";A 4281");		//(= P1_P4_m    P1_P4_datai )) ;4281
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4282");		//(= P1_P4_mf    0b11)) ;4282
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4283");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4283
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4284");		//(= P1_P4_rd    0b1)) ;4284
                                                                P1_P4_m = P1_P4_datai; $display(";A 4285");		//(= P1_P4_m    P1_P4_datai )) ;4285
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4286");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4286
                                                                P1_P4_reg0 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4287");		//(= P1_P4_reg0    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4287
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4288");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4288
                                                                P1_P4_reg1 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4289");		//(= P1_P4_reg1    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4289
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4290");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4290
                                                                P1_P4_reg2 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4291");		//(= P1_P4_reg2    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4291
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4292");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4292
                                                                P1_P4_reg3 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4293");		//(= P1_P4_reg3    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4293
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4294");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4294
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1001 :
                                                begin
                                                    $display(";A 4295");		//(= P1_P4_ff    0b1001)) ;4295
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4296");		//(= P1_P4_mf    0b00)) ;4296
                                                                P1_P4_m = P1_P4_tail; $display(";A 4297");		//(= P1_P4_m    P1_P4_tail )) ;4297
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4298");		//(= P1_P4_mf    0b01)) ;4298
                                                                P1_P4_m = P1_P4_datai; $display(";A 4299");		//(= P1_P4_m    P1_P4_datai )) ;4299
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4300");		//(= P1_P4_addr    P1_P4_tail )) ;4300
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4301");		//(= P1_P4_rd    0b1)) ;4301
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4302");		//(= P1_P4_mf    0b10)) ;4302
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4303");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4303
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4304");		//(= P1_P4_rd    0b1)) ;4304
                                                                P1_P4_m = P1_P4_datai; $display(";A 4305");		//(= P1_P4_m    P1_P4_datai )) ;4305
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4306");		//(= P1_P4_mf    0b11)) ;4306
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4307");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4307
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4308");		//(= P1_P4_rd    0b1)) ;4308
                                                                P1_P4_m = P1_P4_datai; $display(";A 4309");		//(= P1_P4_m    P1_P4_datai )) ;4309
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4310");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4310
                                                                P1_P4_reg0 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4311");		//(= P1_P4_reg0    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4311
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4312");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4312
                                                                P1_P4_reg1 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4313");		//(= P1_P4_reg1    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4313
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4314");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4314
                                                                P1_P4_reg2 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4315");		//(= P1_P4_reg2    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4315
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4316");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4316
                                                                P1_P4_reg3 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4317");		//(= P1_P4_reg3    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4317
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4318");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4318
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1010 :
                                                begin
                                                    $display(";A 4319");		//(= P1_P4_ff    0b1010)) ;4319
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4320");		//(= P1_P4_mf    0b00)) ;4320
                                                                P1_P4_m = P1_P4_tail; $display(";A 4321");		//(= P1_P4_m    P1_P4_tail )) ;4321
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4322");		//(= P1_P4_mf    0b01)) ;4322
                                                                P1_P4_m = P1_P4_datai; $display(";A 4323");		//(= P1_P4_m    P1_P4_datai )) ;4323
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4324");		//(= P1_P4_addr    P1_P4_tail )) ;4324
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4325");		//(= P1_P4_rd    0b1)) ;4325
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4326");		//(= P1_P4_mf    0b10)) ;4326
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4327");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4327
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4328");		//(= P1_P4_rd    0b1)) ;4328
                                                                P1_P4_m = P1_P4_datai; $display(";A 4329");		//(= P1_P4_m    P1_P4_datai )) ;4329
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4330");		//(= P1_P4_mf    0b11)) ;4330
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4331");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4331
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4332");		//(= P1_P4_rd    0b1)) ;4332
                                                                P1_P4_m = P1_P4_datai; $display(";A 4333");		//(= P1_P4_m    P1_P4_datai )) ;4333
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4334");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4334
                                                                P1_P4_reg0 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4335");		//(= P1_P4_reg0    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4335
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4336");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4336
                                                                P1_P4_reg1 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4337");		//(= P1_P4_reg1    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4337
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4338");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4338
                                                                P1_P4_reg2 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4339");		//(= P1_P4_reg2    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4339
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4340");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4340
                                                                P1_P4_reg3 = ((P1_P4_r + P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4341");		//(= P1_P4_reg3    (bv-smod (bv-add P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4341
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4342");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4342
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1011 :
                                                begin
                                                    $display(";A 4343");		//(= P1_P4_ff    0b1011)) ;4343
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4344");		//(= P1_P4_mf    0b00)) ;4344
                                                                P1_P4_m = P1_P4_tail; $display(";A 4345");		//(= P1_P4_m    P1_P4_tail )) ;4345
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4346");		//(= P1_P4_mf    0b01)) ;4346
                                                                P1_P4_m = P1_P4_datai; $display(";A 4347");		//(= P1_P4_m    P1_P4_datai )) ;4347
                                                                P1_P4_addr <= #1 P1_P4_tail; $display(";A 4348");		//(= P1_P4_addr    P1_P4_tail )) ;4348
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4349");		//(= P1_P4_rd    0b1)) ;4349
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4350");		//(= P1_P4_mf    0b10)) ;4350
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 4351");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg1 ) 0b00000000000100000000000000000000))) ;4351
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4352");		//(= P1_P4_rd    0b1)) ;4352
                                                                P1_P4_m = P1_P4_datai; $display(";A 4353");		//(= P1_P4_m    P1_P4_datai )) ;4353
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4354");		//(= P1_P4_mf    0b11)) ;4354
                                                                P1_P4_addr <= #1 ((P1_P4_tail + P1_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 4355");		//(= P1_P4_addr    (bv-smod (bv-add P1_P4_tail  P1_P4_reg2 ) 0b00000000000100000000000000000000))) ;4355
                                                                P1_P4_rd <= #1 1'b1; $display(";A 4356");		//(= P1_P4_rd    0b1)) ;4356
                                                                P1_P4_m = P1_P4_datai; $display(";A 4357");		//(= P1_P4_m    P1_P4_datai )) ;4357
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4358");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4358
                                                                P1_P4_reg0 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4359");		//(= P1_P4_reg0    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4359
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4360");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4360
                                                                P1_P4_reg1 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4361");		//(= P1_P4_reg1    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4361
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4362");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4362
                                                                P1_P4_reg2 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4363");		//(= P1_P4_reg2    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4363
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4364");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4364
                                                                P1_P4_reg3 = ((P1_P4_r - P1_P4_m) % 32'b00000000000000000000000000000000); $display(";A 4365");		//(= P1_P4_reg3    (bv-smod (bv-sub P1_P4_r  P1_P4_m ) 0b00000000000000000000000000000000))) ;4365
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4366");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4366
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1100 :
                                                begin
                                                    $display(";A 4367");		//(= P1_P4_ff    0b1100)) ;4367
                                                    case (P1_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 4368");		//(= P1_P4_mf    0b00)) ;4368
                                                                P1_P4_t = (P1_P4_r / 32'sb00000000000000000000000000000010); $display(";A 4369");		//(= P1_P4_t    (bv-sdiv P1_P4_r  0b00000000000000000000000000000010))) ;4369
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 4370");		//(= P1_P4_mf    0b01)) ;4370
                                                                P1_P4_t = (P1_P4_r / 32'sb00000000000000000000000000000010); $display(";A 4371");		//(= P1_P4_t    (bv-sdiv P1_P4_r  0b00000000000000000000000000000010))) ;4371
                                                                if ((P1_P4_B == 1'b1)) begin
                                                                    $display(";A 4372");		//(= (bv-comp P1_P4_B  0b1)   0b1)) ;4372
                                                                    P1_P4_t = (P1_P4_t % 32'b00100000000000000000000000000000); $display(";A 4374");		//(= P1_P4_t    (bv-smod P1_P4_t  0b00100000000000000000000000000000))) ;4374
                                                                end
                                                                else begin
                                                                    $display(";A 4373");		//(= (bv-comp P1_P4_B  0b1)   0b0)) ;4373
                                                                end
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 4375");		//(= P1_P4_mf    0b10)) ;4375
                                                                P1_P4_t = ((P1_P4_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 4376");		//(= P1_P4_t    (bv-mul (bv-smod P1_P4_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;4376
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 4377");		//(= P1_P4_mf    0b11)) ;4377
                                                                P1_P4_t = ((P1_P4_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 4378");		//(= P1_P4_t    (bv-mul (bv-smod P1_P4_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;4378
                                                                if ((P1_P4_t > 32'b11111111111111111111111111111111)) begin
                                                                    $display(";A 4379");		//(= (bool-to-bv (bv-gt P1_P4_t  0b11111111111111111111111111111111))   0b1)) ;4379
                                                                    P1_P4_B = 1'b1; $display(";A 4381");		//(= P1_P4_B    0b1)) ;4381
                                                                end
                                                                else begin
                                                                    $display(";A 4380");		//(= (bool-to-bv (bv-gt P1_P4_t  0b11111111111111111111111111111111))   0b0)) ;4380
                                                                    P1_P4_B = 1'b0; $display(";A 4382");		//(= P1_P4_B    0b0)) ;4382
                                                                end
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4383");		//(= (and (/= P1_P4_mf  0b00) (/= P1_P4_mf  0b01) (/= P1_P4_mf  0b10) (/= P1_P4_mf  0b11))   true)) ;4383
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                    case (P1_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 4384");		//(= P1_P4_d    0b00000000000000000000000000000000)) ;4384
                                                                P1_P4_reg0 = P1_P4_t; $display(";A 4385");		//(= P1_P4_reg0    P1_P4_t )) ;4385
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 4386");		//(= P1_P4_d    0b00000000000000000000000000000001)) ;4386
                                                                P1_P4_reg1 = P1_P4_t; $display(";A 4387");		//(= P1_P4_reg1    P1_P4_t )) ;4387
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 4388");		//(= P1_P4_d    0b00000000000000000000000000000010)) ;4388
                                                                P1_P4_reg2 = P1_P4_t; $display(";A 4389");		//(= P1_P4_reg2    P1_P4_t )) ;4389
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 4390");		//(= P1_P4_d    0b00000000000000000000000000000011)) ;4390
                                                                P1_P4_reg3 = P1_P4_t; $display(";A 4391");		//(= P1_P4_reg3    P1_P4_t )) ;4391
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 4392");		//(= (and (/= P1_P4_d  0b00000000000000000000000000000000) (/= P1_P4_d  0b00000000000000000000000000000001) (/= P1_P4_d  0b00000000000000000000000000000010) (/= P1_P4_d  0b00000000000000000000000000000011))   true)) ;4392
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1101 :
                                                begin
                                                    $display(";A 4393");		//(= P1_P4_ff    0b1101)) ;4393
                                                    begin
                                                    end
                                                end
                                            4'b1110 :
                                                begin
                                                    $display(";A 4394");		//(= P1_P4_ff    0b1110)) ;4394
                                                    begin
                                                    end
                                                end
                                            4'b1111 :
                                                begin
                                                    $display(";A 4395");		//(= P1_P4_ff    0b1111)) ;4395
                                                    begin
                                                    end
                                                end
                                        endcase
                                    end
                                    else begin
                                        $display(";A 4062");		//(= (bv-not (bv-comp P1_P4_df  0b00000000000000000000000000000111))   0b0)) ;4062
                                        if ((P1_P4_df == 32'b00000000000000000000000000000111)) begin
                                            $display(";A 4396");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000111)   0b1)) ;4396
                                            case (P1_P4_mf)
                                                2'b00 :
                                                    begin
                                                        $display(";A 4398");		//(= P1_P4_mf    0b00)) ;4398
                                                        P1_P4_m = P1_P4_tail; $display(";A 4399");		//(= P1_P4_m    P1_P4_tail )) ;4399
                                                    end
                                                2'b01 :
                                                    begin
                                                        $display(";A 4400");		//(= P1_P4_mf    0b01)) ;4400
                                                        P1_P4_m = P1_P4_tail; $display(";A 4401");		//(= P1_P4_m    P1_P4_tail )) ;4401
                                                    end
                                                2'b10 :
                                                    begin
                                                        $display(";A 4402");		//(= P1_P4_mf    0b10)) ;4402
                                                        P1_P4_m = ((P1_P4_reg1 % 32'b00000000000100000000000000000000) + (P1_P4_tail % 32'b00000000000100000000000000000000)); $display(";A 4403");		//(= P1_P4_m    (bv-add (bv-smod P1_P4_reg1  0b00000000000100000000000000000000) (bv-smod P1_P4_tail  0b00000000000100000000000000000000)))) ;4403
                                                    end
                                                2'b11 :
                                                    begin
                                                        $display(";A 4404");		//(= P1_P4_mf    0b11)) ;4404
                                                        P1_P4_m = ((P1_P4_reg2 % 32'b00000000000100000000000000000000) + (P1_P4_tail % 32'b00000000000100000000000000000000)); $display(";A 4405");		//(= P1_P4_m    (bv-add (bv-smod P1_P4_reg2  0b00000000000100000000000000000000) (bv-smod P1_P4_tail  0b00000000000100000000000000000000)))) ;4405
                                                    end
                                            endcase
                                            P1_P4_addr <= #1 ((P1_P4_m % 32'sb00000000000000000000000000000010) * 32'sb00000000000000000000000000010100); $display(";A 4406");		//(= P1_P4_addr    (bv-mul (bv-smod P1_P4_m  0b00000000000000000000000000000010) 0b00000000000000000000000000010100))) ;4406
                                            P1_P4_wr <= #1 1'b1; $display(";A 4407");		//(= P1_P4_wr    0b1)) ;4407
                                            P1_P4_datao <= #1 P1_P4_r; $display(";A 4408");		//(= P1_P4_datao    P1_P4_r )) ;4408
                                        end
                                        else begin
                                            $display(";A 4397");		//(= (bv-comp P1_P4_df  0b00000000000000000000000000000111)   0b0)) ;4397
                                        end
                                    end
                                end
                        endcase
                        P1_P4_state = 1'sb0; $display(";A 4409");		//(= P1_P4_state    0b0)) ;4409
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6525
    always @(P1_td2 or P1_td1 or P1_din or P1_sel or P1_tad4 or P1_tad3 or P1_ad22 or P1_ad21 or P1_ad12 or P1_ad11 or P1_do4 or P1_do3 or P1_tad1 or P1_ad41 or P1_wr4 or P1_tad2 or P1_ad31 or P1_wr3 or P1_as11 or P1_as21 or P1_as22 or P1_dc2 or P1_mio2 or P1_wr2 or P1_rd4 or P1_do2 or P1_as12 or P1_dc1 or P1_mio1 or P1_wr1 or P1_rd3 or P1_do1) begin
        P1_di3 <= #1 (P1_do1 % 32'b00000000000100000000000000000000); $display(";A 4410");		//(= P1_di3    (bv-smod P1_do1  0b00000000000100000000000000000000))) ;4410
        P1_r12 <= #1 (~((((P1_rd3 & P1_wr1) & P1_mio1) & P1_dc1) & (~P1_as12))); $display(";A 4411");		//(= P1_r12    (bv-not (bv-and (bv-and (bv-and (bv-and P1_rd3  P1_wr1 ) P1_mio1 ) P1_dc1 ) (bv-not P1_as12 ))))) ;4411
        P1_di4 <= #1 P1_do2; $display(";A 4412");		//(= P1_di4    P1_do2 )) ;4412
        P1_r22 <= #1 (~((((P1_rd4 & P1_wr2) & P1_mio2) & P1_dc2) & (~P1_as22))); $display(";A 4413");		//(= P1_r22    (bv-not (bv-and (bv-and (bv-and (bv-and P1_rd4  P1_wr2 ) P1_mio2 ) P1_dc2 ) (bv-not P1_as22 ))))) ;4413
        P1_r11 <= #1 P1_as21; $display(";A 4414");		//(= P1_r11    P1_as21 )) ;4414
        P1_r21 <= #1 P1_as11; $display(";A 4415");		//(= P1_r21    P1_as11 )) ;4415
        if ((P1_wr3 == 1'b1)) begin
            $display(";A 4416");		//(= (bv-comp P1_wr3  0b1)   0b1)) ;4416
            P1_tad3 <= #1 P1_ad31; $display(";A 4418");		//(= P1_tad3    P1_ad31 )) ;4418
        end
        else begin
            $display(";A 4417");		//(= (bv-comp P1_wr3  0b1)   0b0)) ;4417
            P1_tad3 <= #1 (P1_tad2 % 30'b000000000100000000000000000000); $display(";A 4419");		//(= P1_tad3    (bv-smod P1_tad2  0b000000000100000000000000000000))) ;4419
        end
        if ((P1_wr4 == 1'b1)) begin
            $display(";A 4420");		//(= (bv-comp P1_wr4  0b1)   0b1)) ;4420
            P1_tad4 <= #1 P1_ad41; $display(";A 4422");		//(= P1_tad4    P1_ad41 )) ;4422
        end
        else begin
            $display(";A 4421");		//(= (bv-comp P1_wr4  0b1)   0b0)) ;4421
            P1_tad4 <= #1 (P1_tad1 % 30'b000000000100000000000000000000); $display(";A 4423");		//(= P1_tad4    (bv-smod P1_tad1  0b000000000100000000000000000000))) ;4423
        end
        if ((P1_do3 > 32'b00010000000000000000000000000000)) begin
            $display(";A 4424");		//(= (bool-to-bv (bv-gt P1_do3  0b00010000000000000000000000000000))   0b1)) ;4424
            P1_tad1 <= #1 P1_ad11; $display(";A 4426");		//(= P1_tad1    P1_ad11 )) ;4426
        end
        else begin
            $display(";A 4425");		//(= (bool-to-bv (bv-gt P1_do3  0b00010000000000000000000000000000))   0b0)) ;4425
            P1_tad1 <= #1 P1_ad12; $display(";A 4427");		//(= P1_tad1    P1_ad12 )) ;4427
        end
        if ((P1_do4 > 32'b00100000000000000000000000000000)) begin
            $display(";A 4428");		//(= (bool-to-bv (bv-gt P1_do4  0b00100000000000000000000000000000))   0b1)) ;4428
            P1_tad2 <= #1 P1_ad21; $display(";A 4430");		//(= P1_tad2    P1_ad21 )) ;4430
        end
        else begin
            $display(";A 4429");		//(= (bool-to-bv (bv-gt P1_do4  0b00100000000000000000000000000000))   0b0)) ;4429
            P1_tad2 <= #1 P1_ad22; $display(";A 4431");		//(= P1_tad2    P1_ad22 )) ;4431
        end
        P1_dout <= #1 ((P1_tad3 * P1_tad4) % 20'b10000000000000000000); $display(";A 4432");		//(= P1_dout    (bv-smod (bv-mul P1_tad3  P1_tad4 ) 0b10000000000000000000))) ;4432
        if ((P1_sel == 1'b0)) begin
            $display(";A 4433");		//(= (bv-comp P1_sel  0b0)   0b1)) ;4433
            P1_td1 <= #1 32'sb00000000000000000000000000000000; $display(";A 4435");		//(= P1_td1    0b00000000000000000000000000000000)) ;4435
            P1_td2 <= #1 P1_din; $display(";A 4436");		//(= P1_td2    P1_din )) ;4436
        end
        else begin
            $display(";A 4434");		//(= (bv-comp P1_sel  0b0)   0b0)) ;4434
            P1_td1 <= #1 P1_din; $display(";A 4437");		//(= P1_td1    P1_din )) ;4437
            P1_td2 <= #1 32'sb00000000000000000000000000000000; $display(";A 4438");		//(= P1_td2    0b00000000000000000000000000000000)) ;4438
        end
        P1_di1 <= #1 (P1_do4 * P1_td1); $display(";A 4439");		//(= P1_di1    (bv-mul P1_do4  P1_td1 ))) ;4439
        P1_di2 <= #1 (P1_do3 * P1_td2); $display(";A 4440");		//(= P1_di2    (bv-mul P1_do3  P1_td2 ))) ;4440
        P1_aux <= #1 ((P1_tad1 * P1_tad2) % 30'b000000000000000000000000001000); $display(";A 4441");		//(= P1_aux    (bv-smod (bv-mul P1_tad1  P1_tad2 ) 0b000000000000000000000000001000))) ;4441
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6691
    always @(posedge P2_P1_reset or posedge P2_P1_clock) begin
        if ((P2_P1_reset == 1'b1)) begin
            P2_P1_buf1 <= #1 32'sb00000000000000000000000000000000; $display(";A 4444");		//(= P2_P1_buf1    0b00000000000000000000000000000000)) ;4444
            P2_P1_ready11 <= #1 1'b0; $display(";A 4445");		//(= P2_P1_ready11    0b0)) ;4445
            P2_P1_ready12 <= #1 1'b0; $display(";A 4446");		//(= P2_P1_ready12    0b0)) ;4446
        end
        else begin
            if (((((((P2_P1_addr1 > 30'b100000000000000000000000000000) & (P2_P1_ads1 == 1'b0)) & (P2_P1_mio1 == 1'b1)) & (P2_P1_dc1 == 1'b0)) & (P2_P1_wr1 == 1'b1)) & (P2_P1_be1 == 4'b0000))) begin
                $display(";A 4447");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P1_addr1  0b100000000000000000000000000000)) (bv-comp P2_P1_ads1  0b0)) (bv-comp P2_P1_mio1  0b1)) (bv-comp P2_P1_dc1  0b0)) (bv-comp P2_P1_wr1  0b1)) (bv-comp P2_P1_be1  0b0000))   0b1)) ;4447
                P2_P1_buf1 <= #1 P2_P1_do1; $display(";A 4449");		//(= P2_P1_buf1    P2_P1_do1 )) ;4449
                P2_P1_ready11 <= #1 1'b0; $display(";A 4450");		//(= P2_P1_ready11    0b0)) ;4450
                P2_P1_ready12 <= #1 1'b1; $display(";A 4451");		//(= P2_P1_ready12    0b1)) ;4451
            end
            else begin
                $display(";A 4448");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P1_addr1  0b100000000000000000000000000000)) (bv-comp P2_P1_ads1  0b0)) (bv-comp P2_P1_mio1  0b1)) (bv-comp P2_P1_dc1  0b0)) (bv-comp P2_P1_wr1  0b1)) (bv-comp P2_P1_be1  0b0000))   0b0)) ;4448
                if (((((((P2_P1_addr2 > 30'b100000000000000000000000000000) & (P2_P1_ads2 == 1'b0)) & (P2_P1_mio2 == 1'b1)) & (P2_P1_dc2 == 1'b0)) & (P2_P1_wr2 == 1'b1)) & (P2_P1_be2 == 4'b0000))) begin
                    $display(";A 4452");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P1_addr2  0b100000000000000000000000000000)) (bv-comp P2_P1_ads2  0b0)) (bv-comp P2_P1_mio2  0b1)) (bv-comp P2_P1_dc2  0b0)) (bv-comp P2_P1_wr2  0b1)) (bv-comp P2_P1_be2  0b0000))   0b1)) ;4452
                    P2_P1_buf1 <= #1 P2_P1_do2; $display(";A 4454");		//(= P2_P1_buf1    P2_P1_do2 )) ;4454
                    P2_P1_ready11 <= #1 1'b1; $display(";A 4455");		//(= P2_P1_ready11    0b1)) ;4455
                    P2_P1_ready12 <= #1 1'b0; $display(";A 4456");		//(= P2_P1_ready12    0b0)) ;4456
                end
                else begin
                    $display(";A 4453");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P1_addr2  0b100000000000000000000000000000)) (bv-comp P2_P1_ads2  0b0)) (bv-comp P2_P1_mio2  0b1)) (bv-comp P2_P1_dc2  0b0)) (bv-comp P2_P1_wr2  0b1)) (bv-comp P2_P1_be2  0b0000))   0b0)) ;4453
                    P2_P1_ready11 <= #1 1'b1; $display(";A 4457");		//(= P2_P1_ready11    0b1)) ;4457
                    P2_P1_ready12 <= #1 1'b1; $display(";A 4458");		//(= P2_P1_ready12    0b1)) ;4458
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6720
    always @(posedge P2_P1_reset or posedge P2_P1_clock) begin
        if ((P2_P1_reset == 1'b1)) begin
            P2_P1_buf2 <= #1 32'sb00000000000000000000000000000000; $display(";A 4461");		//(= P2_P1_buf2    0b00000000000000000000000000000000)) ;4461
            P2_P1_ready21 <= #1 1'b0; $display(";A 4462");		//(= P2_P1_ready21    0b0)) ;4462
            P2_P1_ready22 <= #1 1'b0; $display(";A 4463");		//(= P2_P1_ready22    0b0)) ;4463
        end
        else begin
            if (((((((P2_P1_addr2 < 30'b100000000000000000000000000000) & (P2_P1_ads2 == 1'b0)) & (P2_P1_mio2 == 1'b1)) & (P2_P1_dc2 == 1'b0)) & (P2_P1_wr2 == 1'b1)) & (P2_P1_be2 == 4'b0000))) begin
                $display(";A 4464");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P2_P1_addr2  0b100000000000000000000000000000)) (bv-comp P2_P1_ads2  0b0)) (bv-comp P2_P1_mio2  0b1)) (bv-comp P2_P1_dc2  0b0)) (bv-comp P2_P1_wr2  0b1)) (bv-comp P2_P1_be2  0b0000))   0b1)) ;4464
                P2_P1_buf2 <= #1 P2_P1_do2; $display(";A 4466");		//(= P2_P1_buf2    P2_P1_do2 )) ;4466
                P2_P1_ready21 <= #1 1'b0; $display(";A 4467");		//(= P2_P1_ready21    0b0)) ;4467
                P2_P1_ready22 <= #1 1'b1; $display(";A 4468");		//(= P2_P1_ready22    0b1)) ;4468
            end
            else begin
                $display(";A 4465");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P2_P1_addr2  0b100000000000000000000000000000)) (bv-comp P2_P1_ads2  0b0)) (bv-comp P2_P1_mio2  0b1)) (bv-comp P2_P1_dc2  0b0)) (bv-comp P2_P1_wr2  0b1)) (bv-comp P2_P1_be2  0b0000))   0b0)) ;4465
                if ((((((P2_P1_ads3 == 1'b0) & (P2_P1_mio3 == 1'b1)) & (P2_P1_dc3 == 1'b0)) & (P2_P1_wr3 == 1'b0)) & (P2_P1_be3 == 4'b0000))) begin
                    $display(";A 4469");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P2_P1_ads3  0b0) (bv-comp P2_P1_mio3  0b1)) (bv-comp P2_P1_dc3  0b0)) (bv-comp P2_P1_wr3  0b0)) (bv-comp P2_P1_be3  0b0000))   0b1)) ;4469
                    P2_P1_ready21 <= #1 1'b1; $display(";A 4471");		//(= P2_P1_ready21    0b1)) ;4471
                    P2_P1_ready22 <= #1 1'b0; $display(";A 4472");		//(= P2_P1_ready22    0b0)) ;4472
                end
                else begin
                    $display(";A 4470");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P2_P1_ads3  0b0) (bv-comp P2_P1_mio3  0b1)) (bv-comp P2_P1_dc3  0b0)) (bv-comp P2_P1_wr3  0b0)) (bv-comp P2_P1_be3  0b0000))   0b0)) ;4470
                    P2_P1_ready21 <= #1 1'b1; $display(";A 4473");		//(= P2_P1_ready21    0b1)) ;4473
                    P2_P1_ready22 <= #1 1'b1; $display(";A 4474");		//(= P2_P1_ready22    0b1)) ;4474
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6748
    always @(P2_P1_datai or P2_P1_buf1 or P2_P1_addr1) begin
        if ((P2_P1_addr1 > 30'b100000000000000000000000000000)) begin
            $display(";A 4475");		//(= (bool-to-bv (bv-gt P2_P1_addr1  0b100000000000000000000000000000))   0b1)) ;4475
            P2_P1_di1 <= #1 P2_P1_buf1; $display(";A 4477");		//(= P2_P1_di1    P2_P1_buf1 )) ;4477
        end
        else begin
            $display(";A 4476");		//(= (bool-to-bv (bv-gt P2_P1_addr1  0b100000000000000000000000000000))   0b0)) ;4476
            P2_P1_di1 <= #1 P2_P1_datai; $display(";A 4478");		//(= P2_P1_di1    P2_P1_datai )) ;4478
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6754
    always @(P2_P1_buf2 or P2_P1_buf1 or P2_P1_addr2) begin
        if ((P2_P1_addr2 > 30'b100000000000000000000000000000)) begin
            $display(";A 4479");		//(= (bool-to-bv (bv-gt P2_P1_addr2  0b100000000000000000000000000000))   0b1)) ;4479
            P2_P1_di2 <= #1 P2_P1_buf1; $display(";A 4481");		//(= P2_P1_di2    P2_P1_buf1 )) ;4481
        end
        else begin
            $display(";A 4480");		//(= (bool-to-bv (bv-gt P2_P1_addr2  0b100000000000000000000000000000))   0b0)) ;4480
            P2_P1_di2 <= #1 P2_P1_buf2; $display(";A 4482");		//(= P2_P1_di2    P2_P1_buf2 )) ;4482
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6760
    always @(P2_P1_do3 or P2_P1_do2 or P2_P1_do1 or P2_P1_addr3 or P2_P1_addr2) begin
        if ((((P2_P1_do1 < 32'b00000000000000000000000000000000) & (P2_P1_do2 < 32'b00000000000000000000000000000000)) & (P2_P1_do3 < 32'b00000000000000000000000000000000))) begin
            $display(";A 4483");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P2_P1_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P2_P1_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P2_P1_do3  0b00000000000000000000000000000000)))   0b1)) ;4483
            P2_P1_address2 <= #1 P2_P1_addr3; $display(";A 4485");		//(= P2_P1_address2    P2_P1_addr3 )) ;4485
        end
        else begin
            $display(";A 4484");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P2_P1_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P2_P1_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P2_P1_do3  0b00000000000000000000000000000000)))   0b0)) ;4484
            P2_P1_address2 <= #1 P2_P1_addr2; $display(";A 4486");		//(= P2_P1_address2    P2_P1_addr2 )) ;4486
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6766
    always @(P2_P1_ready22 or P2_P1_ready21 or P2_P1_ready12 or P2_P1_ready11 or P2_P1_ready2 or P2_P1_ready1 or P2_P1_ads3 or P2_P1_ads1 or P2_P1_mio3 or P2_P1_dc3 or P2_P1_wr3 or P2_P1_addr1 or P2_P1_do3 or P2_P1_buf2) begin
        P2_P1_di3 <= #1 P2_P1_buf2; $display(";A 4487");		//(= P2_P1_di3    P2_P1_buf2 )) ;4487
        P2_P1_datao <= #1 P2_P1_do3; $display(";A 4488");		//(= P2_P1_datao    P2_P1_do3 )) ;4488
        P2_P1_address1 <= #1 P2_P1_addr1; $display(";A 4489");		//(= P2_P1_address1    P2_P1_addr1 )) ;4489
        P2_P1_wr <= #1 P2_P1_wr3; $display(";A 4490");		//(= P2_P1_wr    P2_P1_wr3 )) ;4490
        P2_P1_dc <= #1 P2_P1_dc3; $display(";A 4491");		//(= P2_P1_dc    P2_P1_dc3 )) ;4491
        P2_P1_mio <= #1 P2_P1_mio3; $display(";A 4492");		//(= P2_P1_mio    P2_P1_mio3 )) ;4492
        P2_P1_ast1 <= #1 P2_P1_ads1; $display(";A 4493");		//(= P2_P1_ast1    P2_P1_ads1 )) ;4493
        P2_P1_ast2 <= #1 P2_P1_ads3; $display(";A 4494");		//(= P2_P1_ast2    P2_P1_ads3 )) ;4494
        P2_P1_rdy1 <= #1 (P2_P1_ready11 & P2_P1_ready1); $display(";A 4495");		//(= P2_P1_rdy1    (bv-and P2_P1_ready11  P2_P1_ready1 ))) ;4495
        P2_P1_rdy2 <= #1 (P2_P1_ready12 & P2_P1_ready21); $display(";A 4496");		//(= P2_P1_rdy2    (bv-and P2_P1_ready12  P2_P1_ready21 ))) ;4496
        P2_P1_rdy3 <= #1 (P2_P1_ready22 & P2_P1_ready2); $display(";A 4497");		//(= P2_P1_rdy3    (bv-and P2_P1_ready22  P2_P1_ready2 ))) ;4497
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:6891
    always @(posedge P2_P1_P1_RESET or posedge P2_P1_P1_CLOCK) begin
        if ((P2_P1_P1_RESET == 1'b1)) begin
            $display(";A 4498");		//(= (bv-comp P2_P1_P1_RESET  0b1)   0b1)) ;4498
            P2_P1_P1_BE_n <= #1 4'b0000; $display(";A 4500");		//(= P2_P1_P1_BE_n    0b0000)) ;4500
            P2_P1_P1_Address <= #1 30'sb000000000000000000000000000000; $display(";A 4501");		//(= P2_P1_P1_Address    0b000000000000000000000000000000)) ;4501
            P2_P1_P1_W_R_n <= #1 1'b0; $display(";A 4502");		//(= P2_P1_P1_W_R_n    0b0)) ;4502
            P2_P1_P1_D_C_n <= #1 1'b0; $display(";A 4503");		//(= P2_P1_P1_D_C_n    0b0)) ;4503
            P2_P1_P1_M_IO_n <= #1 1'b0; $display(";A 4504");		//(= P2_P1_P1_M_IO_n    0b0)) ;4504
            P2_P1_P1_ADS_n <= #1 1'b0; $display(";A 4505");		//(= P2_P1_P1_ADS_n    0b0)) ;4505
            P2_P1_P1_State <= #1 3'sb000; $display(";A 4506");		//(= P2_P1_P1_State    0b000)) ;4506
            P2_P1_P1_StateNA <= #1 1'b0; $display(";A 4507");		//(= P2_P1_P1_StateNA    0b0)) ;4507
            P2_P1_P1_StateBS16 <= #1 1'b0; $display(";A 4508");		//(= P2_P1_P1_StateBS16    0b0)) ;4508
            P2_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 4509");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000000)) ;4509
        end
        else begin
            $display(";A 4499");		//(= (bv-comp P2_P1_P1_RESET  0b1)   0b0)) ;4499
            case (P2_P1_P1_State)
                3'b000 :
                    begin
                        $display(";A 4510");		//(= P2_P1_P1_State    0b000)) ;4510
                        P2_P1_P1_D_C_n <= #1 1'b1; $display(";A 4511");		//(= P2_P1_P1_D_C_n    0b1)) ;4511
                        P2_P1_P1_ADS_n <= #1 1'b1; $display(";A 4512");		//(= P2_P1_P1_ADS_n    0b1)) ;4512
                        P2_P1_P1_State <= #1 3'sb001; $display(";A 4513");		//(= P2_P1_P1_State    0b001)) ;4513
                        P2_P1_P1_StateNA <= #1 1'b1; $display(";A 4514");		//(= P2_P1_P1_StateNA    0b1)) ;4514
                        P2_P1_P1_StateBS16 <= #1 1'b1; $display(";A 4515");		//(= P2_P1_P1_StateBS16    0b1)) ;4515
                        P2_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 4516");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;4516
                        P2_P1_P1_State <= #1 3'sb001; $display(";A 4517");		//(= P2_P1_P1_State    0b001)) ;4517
                    end
                3'b001 :
                    begin
                        $display(";A 4518");		//(= P2_P1_P1_State    0b001)) ;4518
                        if ((P2_P1_P1_RequestPending == 1'b1)) begin
                            $display(";A 4519");		//(= (bv-comp P2_P1_P1_RequestPending  0b1)   0b1)) ;4519
                            P2_P1_P1_State <= #1 3'sb010; $display(";A 4521");		//(= P2_P1_P1_State    0b010)) ;4521
                        end
                        else begin
                            $display(";A 4520");		//(= (bv-comp P2_P1_P1_RequestPending  0b1)   0b0)) ;4520
                            if ((P2_P1_P1_HOLD == 1'b1)) begin
                                $display(";A 4522");		//(= (bv-comp P2_P1_P1_HOLD  0b1)   0b1)) ;4522
                                P2_P1_P1_State <= #1 3'sb101; $display(";A 4524");		//(= P2_P1_P1_State    0b101)) ;4524
                            end
                            else begin
                                $display(";A 4523");		//(= (bv-comp P2_P1_P1_HOLD  0b1)   0b0)) ;4523
                                P2_P1_P1_State <= #1 3'sb001; $display(";A 4525");		//(= P2_P1_P1_State    0b001)) ;4525
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 4526");		//(= P2_P1_P1_State    0b010)) ;4526
                        P2_P1_P1_Address <= #1 ((P2_P1_P1_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 4527");		//(= P2_P1_P1_Address    (bv-smod (bv-sdiv P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;4527
                        P2_P1_P1_BE_n <= #1 P2_P1_P1_ByteEnable; $display(";A 4528");		//(= P2_P1_P1_BE_n    P2_P1_P1_ByteEnable )) ;4528
                        P2_P1_P1_M_IO_n <= #1 P2_P1_P1_MemoryFetch; $display(";A 4529");		//(= P2_P1_P1_M_IO_n    P2_P1_P1_MemoryFetch )) ;4529
                        if ((P2_P1_P1_ReadRequest == 1'b1)) begin
                            $display(";A 4530");		//(= (bv-comp P2_P1_P1_ReadRequest  0b1)   0b1)) ;4530
                            P2_P1_P1_W_R_n <= #1 1'b0; $display(";A 4532");		//(= P2_P1_P1_W_R_n    0b0)) ;4532
                        end
                        else begin
                            $display(";A 4531");		//(= (bv-comp P2_P1_P1_ReadRequest  0b1)   0b0)) ;4531
                            P2_P1_P1_W_R_n <= #1 1'b1; $display(";A 4533");		//(= P2_P1_P1_W_R_n    0b1)) ;4533
                        end
                        if ((P2_P1_P1_CodeFetch == 1'b1)) begin
                            $display(";A 4534");		//(= (bv-comp P2_P1_P1_CodeFetch  0b1)   0b1)) ;4534
                            P2_P1_P1_D_C_n <= #1 1'b0; $display(";A 4536");		//(= P2_P1_P1_D_C_n    0b0)) ;4536
                        end
                        else begin
                            $display(";A 4535");		//(= (bv-comp P2_P1_P1_CodeFetch  0b1)   0b0)) ;4535
                            P2_P1_P1_D_C_n <= #1 1'b1; $display(";A 4537");		//(= P2_P1_P1_D_C_n    0b1)) ;4537
                        end
                        P2_P1_P1_ADS_n <= #1 1'b0; $display(";A 4538");		//(= P2_P1_P1_ADS_n    0b0)) ;4538
                        P2_P1_P1_State <= #1 3'sb011; $display(";A 4539");		//(= P2_P1_P1_State    0b011)) ;4539
                    end
                3'b011 :
                    begin
                        $display(";A 4540");		//(= P2_P1_P1_State    0b011)) ;4540
                        if ((((P2_P1_P1_READY_n == 1'b0) & (P2_P1_P1_HOLD == 1'b0)) & (P2_P1_P1_RequestPending == 1'b1))) begin
                            $display(";A 4541");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b1))   0b1)) ;4541
                            P2_P1_P1_State <= #1 3'sb010; $display(";A 4543");		//(= P2_P1_P1_State    0b010)) ;4543
                        end
                        else begin
                            $display(";A 4542");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b1))   0b0)) ;4542
                            if (((P2_P1_P1_READY_n == 1'b1) & (P2_P1_P1_NA_n == 1'b1))) begin
                                $display(";A 4544");		//(= (bv-and (bv-comp P2_P1_P1_READY_n  0b1) (bv-comp P2_P1_P1_NA_n  0b1))   0b1)) ;4544
                            end
                            else begin
                                $display(";A 4545");		//(= (bv-and (bv-comp P2_P1_P1_READY_n  0b1) (bv-comp P2_P1_P1_NA_n  0b1))   0b0)) ;4545
                                if ((((P2_P1_P1_RequestPending == 1'b1) | (P2_P1_P1_HOLD == 1'b1)) & ((P2_P1_P1_READY_n == 1'b1) & (P2_P1_P1_NA_n == 1'b0)))) begin
                                    $display(";A 4546");		//(= (bv-and (bv-or (bv-comp P2_P1_P1_RequestPending  0b1) (bv-comp P2_P1_P1_HOLD  0b1)) (bv-and (bv-comp P2_P1_P1_READY_n  0b1) (bv-comp P2_P1_P1_NA_n  0b0)))   0b1)) ;4546
                                    P2_P1_P1_State <= #1 3'sb111; $display(";A 4548");		//(= P2_P1_P1_State    0b111)) ;4548
                                end
                                else begin
                                    $display(";A 4547");		//(= (bv-and (bv-or (bv-comp P2_P1_P1_RequestPending  0b1) (bv-comp P2_P1_P1_HOLD  0b1)) (bv-and (bv-comp P2_P1_P1_READY_n  0b1) (bv-comp P2_P1_P1_NA_n  0b0)))   0b0)) ;4547
                                    if (((((P2_P1_P1_RequestPending == 1'b1) & (P2_P1_P1_HOLD == 1'b0)) & (P2_P1_P1_READY_n == 1'b1)) & (P2_P1_P1_NA_n == 1'b0))) begin
                                        $display(";A 4549");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P1_P1_RequestPending  0b1) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_READY_n  0b1)) (bv-comp P2_P1_P1_NA_n  0b0))   0b1)) ;4549
                                        P2_P1_P1_State <= #1 3'sb110; $display(";A 4551");		//(= P2_P1_P1_State    0b110)) ;4551
                                    end
                                    else begin
                                        $display(";A 4550");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P1_P1_RequestPending  0b1) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_READY_n  0b1)) (bv-comp P2_P1_P1_NA_n  0b0))   0b0)) ;4550
                                        if ((((P2_P1_P1_RequestPending == 1'b0) & (P2_P1_P1_HOLD == 1'b0)) & (P2_P1_P1_READY_n == 1'b0))) begin
                                            $display(";A 4552");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_RequestPending  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_READY_n  0b0))   0b1)) ;4552
                                            P2_P1_P1_State <= #1 3'sb001; $display(";A 4554");		//(= P2_P1_P1_State    0b001)) ;4554
                                        end
                                        else begin
                                            $display(";A 4553");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_RequestPending  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_READY_n  0b0))   0b0)) ;4553
                                            if (((P2_P1_P1_HOLD == 1'b1) & (P2_P1_P1_READY_n == 1'b1))) begin
                                                $display(";A 4555");		//(= (bv-and (bv-comp P2_P1_P1_HOLD  0b1) (bv-comp P2_P1_P1_READY_n  0b1))   0b1)) ;4555
                                                P2_P1_P1_State <= #1 3'sb101; $display(";A 4557");		//(= P2_P1_P1_State    0b101)) ;4557
                                            end
                                            else begin
                                                $display(";A 4556");		//(= (bv-and (bv-comp P2_P1_P1_HOLD  0b1) (bv-comp P2_P1_P1_READY_n  0b1))   0b0)) ;4556
                                                P2_P1_P1_State <= #1 3'sb011; $display(";A 4558");		//(= P2_P1_P1_State    0b011)) ;4558
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P2_P1_P1_StateBS16 <= #1 P2_P1_P1_BS16_n; $display(";A 4559");		//(= P2_P1_P1_StateBS16    P2_P1_P1_BS16_n )) ;4559
                        if ((P2_P1_P1_BS16_n == 1'b0)) begin
                            $display(";A 4560");		//(= (bv-comp P2_P1_P1_BS16_n  0b0)   0b1)) ;4560
                            P2_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 4562");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000001)) ;4562
                        end
                        else begin
                            $display(";A 4561");		//(= (bv-comp P2_P1_P1_BS16_n  0b0)   0b0)) ;4561
                            P2_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 4563");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;4563
                        end
                        P2_P1_P1_StateNA <= #1 P2_P1_P1_NA_n; $display(";A 4564");		//(= P2_P1_P1_StateNA    P2_P1_P1_NA_n )) ;4564
                        P2_P1_P1_ADS_n <= #1 1'b1; $display(";A 4565");		//(= P2_P1_P1_ADS_n    0b1)) ;4565
                    end
                3'b100 :
                    begin
                        $display(";A 4566");		//(= P2_P1_P1_State    0b100)) ;4566
                        if ((((P2_P1_P1_NA_n == 1'b0) & (P2_P1_P1_HOLD == 1'b0)) & (P2_P1_P1_RequestPending == 1'b1))) begin
                            $display(";A 4567");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_NA_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b1))   0b1)) ;4567
                            P2_P1_P1_State <= #1 3'sb110; $display(";A 4569");		//(= P2_P1_P1_State    0b110)) ;4569
                        end
                        else begin
                            $display(";A 4568");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_NA_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b1))   0b0)) ;4568
                            if (((P2_P1_P1_NA_n == 1'b0) & ((P2_P1_P1_HOLD == 1'b1) | (P2_P1_P1_RequestPending == 1'b0)))) begin
                                $display(";A 4570");		//(= (bv-and (bv-comp P2_P1_P1_NA_n  0b0) (bv-or (bv-comp P2_P1_P1_HOLD  0b1) (bv-comp P2_P1_P1_RequestPending  0b0)))   0b1)) ;4570
                                P2_P1_P1_State <= #1 3'sb111; $display(";A 4572");		//(= P2_P1_P1_State    0b111)) ;4572
                            end
                            else begin
                                $display(";A 4571");		//(= (bv-and (bv-comp P2_P1_P1_NA_n  0b0) (bv-or (bv-comp P2_P1_P1_HOLD  0b1) (bv-comp P2_P1_P1_RequestPending  0b0)))   0b0)) ;4571
                                if ((P2_P1_P1_NA_n == 1'b1)) begin
                                    $display(";A 4573");		//(= (bv-comp P2_P1_P1_NA_n  0b1)   0b1)) ;4573
                                    P2_P1_P1_State <= #1 3'sb011; $display(";A 4575");		//(= P2_P1_P1_State    0b011)) ;4575
                                end
                                else begin
                                    $display(";A 4574");		//(= (bv-comp P2_P1_P1_NA_n  0b1)   0b0)) ;4574
                                    P2_P1_P1_State <= #1 3'sb100; $display(";A 4576");		//(= P2_P1_P1_State    0b100)) ;4576
                                end
                            end
                        end
                        P2_P1_P1_StateBS16 <= #1 P2_P1_P1_BS16_n; $display(";A 4577");		//(= P2_P1_P1_StateBS16    P2_P1_P1_BS16_n )) ;4577
                        if ((P2_P1_P1_BS16_n == 1'b0)) begin
                            $display(";A 4578");		//(= (bv-comp P2_P1_P1_BS16_n  0b0)   0b1)) ;4578
                            P2_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 4580");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000001)) ;4580
                        end
                        else begin
                            $display(";A 4579");		//(= (bv-comp P2_P1_P1_BS16_n  0b0)   0b0)) ;4579
                            P2_P1_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 4581");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;4581
                        end
                        P2_P1_P1_StateNA <= #1 P2_P1_P1_NA_n; $display(";A 4582");		//(= P2_P1_P1_StateNA    P2_P1_P1_NA_n )) ;4582
                        P2_P1_P1_ADS_n <= #1 1'b1; $display(";A 4583");		//(= P2_P1_P1_ADS_n    0b1)) ;4583
                    end
                3'b101 :
                    begin
                        $display(";A 4584");		//(= P2_P1_P1_State    0b101)) ;4584
                        if (((P2_P1_P1_HOLD == 1'b0) & (P2_P1_P1_RequestPending == 1'b1))) begin
                            $display(";A 4585");		//(= (bv-and (bv-comp P2_P1_P1_HOLD  0b0) (bv-comp P2_P1_P1_RequestPending  0b1))   0b1)) ;4585
                            P2_P1_P1_State <= #1 3'sb010; $display(";A 4587");		//(= P2_P1_P1_State    0b010)) ;4587
                        end
                        else begin
                            $display(";A 4586");		//(= (bv-and (bv-comp P2_P1_P1_HOLD  0b0) (bv-comp P2_P1_P1_RequestPending  0b1))   0b0)) ;4586
                            if (((P2_P1_P1_HOLD == 1'b0) & (P2_P1_P1_RequestPending == 1'b0))) begin
                                $display(";A 4588");		//(= (bv-and (bv-comp P2_P1_P1_HOLD  0b0) (bv-comp P2_P1_P1_RequestPending  0b0))   0b1)) ;4588
                                P2_P1_P1_State <= #1 3'sb001; $display(";A 4590");		//(= P2_P1_P1_State    0b001)) ;4590
                            end
                            else begin
                                $display(";A 4589");		//(= (bv-and (bv-comp P2_P1_P1_HOLD  0b0) (bv-comp P2_P1_P1_RequestPending  0b0))   0b0)) ;4589
                                P2_P1_P1_State <= #1 3'sb101; $display(";A 4591");		//(= P2_P1_P1_State    0b101)) ;4591
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 4592");		//(= P2_P1_P1_State    0b110)) ;4592
                        P2_P1_P1_Address <= #1 ((P2_P1_P1_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 4593");		//(= P2_P1_P1_Address    (bv-smod (bv-sdiv P2_P1_P1_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;4593
                        P2_P1_P1_BE_n <= #1 P2_P1_P1_ByteEnable; $display(";A 4594");		//(= P2_P1_P1_BE_n    P2_P1_P1_ByteEnable )) ;4594
                        P2_P1_P1_M_IO_n <= #1 P2_P1_P1_MemoryFetch; $display(";A 4595");		//(= P2_P1_P1_M_IO_n    P2_P1_P1_MemoryFetch )) ;4595
                        if ((P2_P1_P1_ReadRequest == 1'b1)) begin
                            $display(";A 4596");		//(= (bv-comp P2_P1_P1_ReadRequest  0b1)   0b1)) ;4596
                            P2_P1_P1_W_R_n <= #1 1'b0; $display(";A 4598");		//(= P2_P1_P1_W_R_n    0b0)) ;4598
                        end
                        else begin
                            $display(";A 4597");		//(= (bv-comp P2_P1_P1_ReadRequest  0b1)   0b0)) ;4597
                            P2_P1_P1_W_R_n <= #1 1'b1; $display(";A 4599");		//(= P2_P1_P1_W_R_n    0b1)) ;4599
                        end
                        if ((P2_P1_P1_CodeFetch == 1'b1)) begin
                            $display(";A 4600");		//(= (bv-comp P2_P1_P1_CodeFetch  0b1)   0b1)) ;4600
                            P2_P1_P1_D_C_n <= #1 1'b0; $display(";A 4602");		//(= P2_P1_P1_D_C_n    0b0)) ;4602
                        end
                        else begin
                            $display(";A 4601");		//(= (bv-comp P2_P1_P1_CodeFetch  0b1)   0b0)) ;4601
                            P2_P1_P1_D_C_n <= #1 1'b1; $display(";A 4603");		//(= P2_P1_P1_D_C_n    0b1)) ;4603
                        end
                        P2_P1_P1_ADS_n <= #1 1'b0; $display(";A 4604");		//(= P2_P1_P1_ADS_n    0b0)) ;4604
                        if ((P2_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 4605");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4605
                            P2_P1_P1_State <= #1 3'sb100; $display(";A 4607");		//(= P2_P1_P1_State    0b100)) ;4607
                        end
                        else begin
                            $display(";A 4606");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4606
                            P2_P1_P1_State <= #1 3'sb110; $display(";A 4608");		//(= P2_P1_P1_State    0b110)) ;4608
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 4609");		//(= P2_P1_P1_State    0b111)) ;4609
                        if ((((P2_P1_P1_READY_n == 1'b1) & (P2_P1_P1_RequestPending == 1'b1)) & (P2_P1_P1_HOLD == 1'b0))) begin
                            $display(";A 4610");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b1) (bv-comp P2_P1_P1_RequestPending  0b1)) (bv-comp P2_P1_P1_HOLD  0b0))   0b1)) ;4610
                            P2_P1_P1_State <= #1 3'sb110; $display(";A 4612");		//(= P2_P1_P1_State    0b110)) ;4612
                        end
                        else begin
                            $display(";A 4611");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b1) (bv-comp P2_P1_P1_RequestPending  0b1)) (bv-comp P2_P1_P1_HOLD  0b0))   0b0)) ;4611
                            if (((P2_P1_P1_READY_n == 1'b0) & (P2_P1_P1_HOLD == 1'b1))) begin
                                $display(";A 4613");		//(= (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b1))   0b1)) ;4613
                                P2_P1_P1_State <= #1 3'sb101; $display(";A 4615");		//(= P2_P1_P1_State    0b101)) ;4615
                            end
                            else begin
                                $display(";A 4614");		//(= (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b1))   0b0)) ;4614
                                if ((((P2_P1_P1_READY_n == 1'b0) & (P2_P1_P1_HOLD == 1'b0)) & (P2_P1_P1_RequestPending == 1'b1))) begin
                                    $display(";A 4616");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b1))   0b1)) ;4616
                                    P2_P1_P1_State <= #1 3'sb010; $display(";A 4618");		//(= P2_P1_P1_State    0b010)) ;4618
                                end
                                else begin
                                    $display(";A 4617");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b1))   0b0)) ;4617
                                    if ((((P2_P1_P1_READY_n == 1'b0) & (P2_P1_P1_HOLD == 1'b0)) & (P2_P1_P1_RequestPending == 1'b0))) begin
                                        $display(";A 4619");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b0))   0b1)) ;4619
                                        P2_P1_P1_State <= #1 3'sb001; $display(";A 4621");		//(= P2_P1_P1_State    0b001)) ;4621
                                    end
                                    else begin
                                        $display(";A 4620");		//(= (bv-and (bv-and (bv-comp P2_P1_P1_READY_n  0b0) (bv-comp P2_P1_P1_HOLD  0b0)) (bv-comp P2_P1_P1_RequestPending  0b0))   0b0)) ;4620
                                        P2_P1_P1_State <= #1 3'sb111; $display(";A 4622");		//(= P2_P1_P1_State    0b111)) ;4622
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:7035
    always @(posedge P2_P1_P1_RESET or posedge P2_P1_P1_CLOCK) begin
        if ((P2_P1_P1_RESET == 1'b1)) begin
            $display(";A 4623");		//(= (bv-comp P2_P1_P1_RESET  0b1)   0b1)) ;4623
            P2_P1_P1_State2 = 4'sb0000; $display(";A 4625");		//(= P2_P1_P1_State2    0b0000)) ;4625
            P2_P1_P1_InstQueue[0] = 8'b00000000; $display(";A 4626");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4626
            P2_P1_P1_InstQueue[1] = 8'b00000000; $display(";A 4627");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4627
            P2_P1_P1_InstQueue[2] = 8'b00000000; $display(";A 4628");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4628
            P2_P1_P1_InstQueue[3] = 8'b00000000; $display(";A 4629");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4629
            P2_P1_P1_InstQueue[4] = 8'b00000000; $display(";A 4630");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4630
            P2_P1_P1_InstQueue[5] = 8'b00000000; $display(";A 4631");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4631
            P2_P1_P1_InstQueue[6] = 8'b00000000; $display(";A 4632");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4632
            P2_P1_P1_InstQueue[7] = 8'b00000000; $display(";A 4633");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4633
            P2_P1_P1_InstQueue[8] = 8'b00000000; $display(";A 4634");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4634
            P2_P1_P1_InstQueue[9] = 8'b00000000; $display(";A 4635");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4635
            P2_P1_P1_InstQueue[10] = 8'b00000000; $display(";A 4636");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4636
            P2_P1_P1_InstQueue[11] = 8'b00000000; $display(";A 4637");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4637
            P2_P1_P1_InstQueue[12] = 8'b00000000; $display(";A 4638");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4638
            P2_P1_P1_InstQueue[13] = 8'b00000000; $display(";A 4639");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4639
            P2_P1_P1_InstQueue[14] = 8'b00000000; $display(";A 4640");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4640
            P2_P1_P1_InstQueue[15] = 8'b00000000; $display(";A 4641");		//(= P2_P1_P1_InstQueue    0b00000000)) ;4641
            P2_P1_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 4642");		//(= P2_P1_P1_InstQueueRd_Addr    0b00000)) ;4642
            P2_P1_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 4643");		//(= P2_P1_P1_InstQueueWr_Addr    0b00000)) ;4643
            P2_P1_P1_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 4644");		//(= P2_P1_P1_InstAddrPointer    0b00000000000000000000000000000000)) ;4644
            P2_P1_P1_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 4645");		//(= P2_P1_P1_PhyAddrPointer    0b00000000000000000000000000000000)) ;4645
            P2_P1_P1_Extended = 1'b0; $display(";A 4646");		//(= P2_P1_P1_Extended    0b0)) ;4646
            P2_P1_P1_More = 1'b0; $display(";A 4647");		//(= P2_P1_P1_More    0b0)) ;4647
            P2_P1_P1_Flush = 1'b0; $display(";A 4648");		//(= P2_P1_P1_Flush    0b0)) ;4648
            P2_P1_P1_lWord = 16'sb0000000000000000; $display(";A 4649");		//(= P2_P1_P1_lWord    0b0000000000000000)) ;4649
            P2_P1_P1_uWord = 15'sb000000000000000; $display(";A 4650");		//(= P2_P1_P1_uWord    0b000000000000000)) ;4650
            P2_P1_P1_fWord = 32'sb00000000000000000000000000000000; $display(";A 4651");		//(= P2_P1_P1_fWord    0b00000000000000000000000000000000)) ;4651
            P2_P1_P1_CodeFetch <= #1 1'b0; $display(";A 4652");		//(= P2_P1_P1_CodeFetch    0b0)) ;4652
            P2_P1_P1_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 4653");		//(= P2_P1_P1_Datao    0b00000000000000000000000000000000)) ;4653
            P2_P1_P1_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 4654");		//(= P2_P1_P1_EAX    0b00000000000000000000000000000000)) ;4654
            P2_P1_P1_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 4655");		//(= P2_P1_P1_EBX    0b00000000000000000000000000000000)) ;4655
            P2_P1_P1_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 4656");		//(= P2_P1_P1_rEIP    0b00000000000000000000000000000000)) ;4656
            P2_P1_P1_ReadRequest <= #1 1'b0; $display(";A 4657");		//(= P2_P1_P1_ReadRequest    0b0)) ;4657
            P2_P1_P1_MemoryFetch <= #1 1'b0; $display(";A 4658");		//(= P2_P1_P1_MemoryFetch    0b0)) ;4658
            P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4659");		//(= P2_P1_P1_RequestPending    0b0)) ;4659
        end
        else begin
            $display(";A 4624");		//(= (bv-comp P2_P1_P1_RESET  0b1)   0b0)) ;4624
            case (P2_P1_P1_State2)
                4'b0000 :
                    begin
                        $display(";A 4660");		//(= P2_P1_P1_State2    0b0000)) ;4660
                        P2_P1_P1_PhyAddrPointer = P2_P1_P1_rEIP; $display(";A 4661");		//(= P2_P1_P1_PhyAddrPointer    P2_P1_P1_rEIP )) ;4661
                        P2_P1_P1_InstAddrPointer = P2_P1_P1_PhyAddrPointer; $display(";A 4662");		//(= P2_P1_P1_InstAddrPointer    P2_P1_P1_PhyAddrPointer )) ;4662
                        P2_P1_P1_State2 = 4'sb0001; $display(";A 4663");		//(= P2_P1_P1_State2    0b0001)) ;4663
                        P2_P1_P1_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 4664");		//(= P2_P1_P1_rEIP    0b00000000000011111111111111110000)) ;4664
                        P2_P1_P1_ReadRequest <= #1 1'b1; $display(";A 4665");		//(= P2_P1_P1_ReadRequest    0b1)) ;4665
                        P2_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 4666");		//(= P2_P1_P1_MemoryFetch    0b1)) ;4666
                        P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4667");		//(= P2_P1_P1_RequestPending    0b1)) ;4667
                    end
                4'b0001 :
                    begin
                        $display(";A 4668");		//(= P2_P1_P1_State2    0b0001)) ;4668
                        P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4669");		//(= P2_P1_P1_RequestPending    0b1)) ;4669
                        P2_P1_P1_ReadRequest <= #1 1'b1; $display(";A 4670");		//(= P2_P1_P1_ReadRequest    0b1)) ;4670
                        P2_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 4671");		//(= P2_P1_P1_MemoryFetch    0b1)) ;4671
                        P2_P1_P1_CodeFetch <= #1 1'b1; $display(";A 4672");		//(= P2_P1_P1_CodeFetch    0b1)) ;4672
                        if ((P2_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 4673");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4673
                            P2_P1_P1_State2 = 4'sb0010; $display(";A 4675");		//(= P2_P1_P1_State2    0b0010)) ;4675
                        end
                        else begin
                            $display(";A 4674");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4674
                            P2_P1_P1_State2 = 4'sb0001; $display(";A 4676");		//(= P2_P1_P1_State2    0b0001)) ;4676
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 4677");		//(= P2_P1_P1_State2    0b0010)) ;4677
                        P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4678");		//(= P2_P1_P1_RequestPending    0b0)) ;4678
                        P2_P1_P1_InstQueue[P2_P1_P1_InstQueueWr_Addr] = (P2_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 4679");		//(= P2_P1_P1_InstQueue    (bv-smod P2_P1_P1_Datai  0b00000000000000000000000100000000))) ;4679
                        P2_P1_P1_InstQueueWr_Addr = ((P2_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4680");		//(= P2_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4680
                        P2_P1_P1_InstQueue[P2_P1_P1_InstQueueWr_Addr] = (P2_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 4681");		//(= P2_P1_P1_InstQueue    (bv-smod P2_P1_P1_Datai  0b00000000000000000000000100000000))) ;4681
                        P2_P1_P1_InstQueueWr_Addr = ((P2_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4682");		//(= P2_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4682
                        if ((P2_P1_P1_StateBS16 == 1'b1)) begin
                            $display(";A 4683");		//(= (bv-comp P2_P1_P1_StateBS16  0b1)   0b1)) ;4683
                            P2_P1_P1_InstQueue[P2_P1_P1_InstQueueWr_Addr] = ((P2_P1_P1_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 4685");		//(= P2_P1_P1_InstQueue    (bv-smod (bv-sdiv P2_P1_P1_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;4685
                            P2_P1_P1_InstQueueWr_Addr = ((P2_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4686");		//(= P2_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4686
                            P2_P1_P1_InstQueue[P2_P1_P1_InstQueueWr_Addr] = ((P2_P1_P1_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 4687");		//(= P2_P1_P1_InstQueue    (bv-smod (bv-sdiv P2_P1_P1_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;4687
                            P2_P1_P1_InstQueueWr_Addr = ((P2_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4688");		//(= P2_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4688
                            P2_P1_P1_PhyAddrPointer = (P2_P1_P1_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 4689");		//(= P2_P1_P1_PhyAddrPointer    (bv-add P2_P1_P1_PhyAddrPointer  0b00000000000000000000000000000100))) ;4689
                            P2_P1_P1_State2 = 4'sb0101; $display(";A 4690");		//(= P2_P1_P1_State2    0b0101)) ;4690
                        end
                        else begin
                            $display(";A 4684");		//(= (bv-comp P2_P1_P1_StateBS16  0b1)   0b0)) ;4684
                            P2_P1_P1_PhyAddrPointer = (P2_P1_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4691");		//(= P2_P1_P1_PhyAddrPointer    (bv-add P2_P1_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;4691
                            if ((P2_P1_P1_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 4692");		//(= (bool-to-bv (bv-slt P2_P1_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;4692
                                P2_P1_P1_rEIP <= #1 (-P2_P1_P1_PhyAddrPointer); $display(";A 4694");		//(= P2_P1_P1_rEIP    (bv-neg P2_P1_P1_PhyAddrPointer ))) ;4694
                            end
                            else begin
                                $display(";A 4693");		//(= (bool-to-bv (bv-slt P2_P1_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;4693
                                P2_P1_P1_rEIP <= #1 P2_P1_P1_PhyAddrPointer; $display(";A 4695");		//(= P2_P1_P1_rEIP    P2_P1_P1_PhyAddrPointer )) ;4695
                            end
                            P2_P1_P1_State2 = 4'sb0011; $display(";A 4696");		//(= P2_P1_P1_State2    0b0011)) ;4696
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 4697");		//(= P2_P1_P1_State2    0b0011)) ;4697
                        P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4698");		//(= P2_P1_P1_RequestPending    0b1)) ;4698
                        if ((P2_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 4699");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4699
                            P2_P1_P1_State2 = 4'sb0100; $display(";A 4701");		//(= P2_P1_P1_State2    0b0100)) ;4701
                        end
                        else begin
                            $display(";A 4700");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4700
                            P2_P1_P1_State2 = 4'sb0011; $display(";A 4702");		//(= P2_P1_P1_State2    0b0011)) ;4702
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 4703");		//(= P2_P1_P1_State2    0b0100)) ;4703
                        P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4704");		//(= P2_P1_P1_RequestPending    0b0)) ;4704
                        P2_P1_P1_InstQueue[P2_P1_P1_InstQueueWr_Addr] = (P2_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 4705");		//(= P2_P1_P1_InstQueue    (bv-smod P2_P1_P1_Datai  0b00000000000000000000000100000000))) ;4705
                        P2_P1_P1_InstQueueWr_Addr = ((P2_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4706");		//(= P2_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4706
                        P2_P1_P1_InstQueue[P2_P1_P1_InstQueueWr_Addr] = (P2_P1_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 4707");		//(= P2_P1_P1_InstQueue    (bv-smod P2_P1_P1_Datai  0b00000000000000000000000100000000))) ;4707
                        P2_P1_P1_InstQueueWr_Addr = ((P2_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4708");		//(= P2_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4708
                        P2_P1_P1_PhyAddrPointer = (P2_P1_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4709");		//(= P2_P1_P1_PhyAddrPointer    (bv-add P2_P1_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;4709
                        P2_P1_P1_State2 = 4'sb0101; $display(";A 4710");		//(= P2_P1_P1_State2    0b0101)) ;4710
                    end
                4'b0101 :
                    begin
                        $display(";A 4711");		//(= P2_P1_P1_State2    0b0101)) ;4711
                        case (P2_P1_P1_InstQueue[P2_P1_P1_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 4712");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b10010000)) ;4712
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4713");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4713
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4714");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4714
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4715");		//(= P2_P1_P1_Flush    0b0)) ;4715
                                    P2_P1_P1_More = 1'b0; $display(";A 4716");		//(= P2_P1_P1_More    0b0)) ;4716
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 4717");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b01100110)) ;4717
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4718");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4718
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4719");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4719
                                    P2_P1_P1_Extended = 1'b1; $display(";A 4720");		//(= P2_P1_P1_Extended    0b1)) ;4720
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4721");		//(= P2_P1_P1_Flush    0b0)) ;4721
                                    P2_P1_P1_More = 1'b0; $display(";A 4722");		//(= P2_P1_P1_More    0b0)) ;4722
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 4723");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b11101011)) ;4723
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 4724");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;4724
                                        if ((P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 4726");		//(= (bool-to-bv (bv-gt P2_P1_P1_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;4726
                                            P2_P1_P1_PhyAddrPointer = ((P2_P1_P1_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 4728");		//(= P2_P1_P1_PhyAddrPointer    (bv-sub (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P2_P1_P1_InstQueue 0 )))) ;4728
                                            P2_P1_P1_InstAddrPointer = P2_P1_P1_PhyAddrPointer; $display(";A 4729");		//(= P2_P1_P1_InstAddrPointer    P2_P1_P1_PhyAddrPointer )) ;4729
                                        end
                                        else begin
                                            $display(";A 4727");		//(= (bool-to-bv (bv-gt P2_P1_P1_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;4727
                                            P2_P1_P1_PhyAddrPointer = ((P2_P1_P1_InstAddrPointer + 32'b00000000000000000000000000000010) + P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 4730");		//(= P2_P1_P1_PhyAddrPointer    (bv-add (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000010) P2_P1_P1_InstQueue 0 ))) ;4730
                                            P2_P1_P1_InstAddrPointer = P2_P1_P1_PhyAddrPointer; $display(";A 4731");		//(= P2_P1_P1_InstAddrPointer    P2_P1_P1_PhyAddrPointer )) ;4731
                                        end
                                        P2_P1_P1_Flush = 1'b1; $display(";A 4732");		//(= P2_P1_P1_Flush    0b1)) ;4732
                                        P2_P1_P1_More = 1'b0; $display(";A 4733");		//(= P2_P1_P1_More    0b0)) ;4733
                                    end
                                    else begin
                                        $display(";A 4725");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;4725
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4734");		//(= P2_P1_P1_Flush    0b0)) ;4734
                                        P2_P1_P1_More = 1'b1; $display(";A 4735");		//(= P2_P1_P1_More    0b1)) ;4735
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 4736");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b11101001)) ;4736
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 4737");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;4737
                                        P2_P1_P1_PhyAddrPointer = ((P2_P1_P1_InstAddrPointer + 32'b00000000000000000000000000000101) + P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 4739");		//(= P2_P1_P1_PhyAddrPointer    (bv-add (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000101) P2_P1_P1_InstQueue 0 ))) ;4739
                                        P2_P1_P1_InstAddrPointer = P2_P1_P1_PhyAddrPointer; $display(";A 4740");		//(= P2_P1_P1_InstAddrPointer    P2_P1_P1_PhyAddrPointer )) ;4740
                                        P2_P1_P1_Flush = 1'b1; $display(";A 4741");		//(= P2_P1_P1_Flush    0b1)) ;4741
                                        P2_P1_P1_More = 1'b0; $display(";A 4742");		//(= P2_P1_P1_More    0b0)) ;4742
                                    end
                                    else begin
                                        $display(";A 4738");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;4738
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4743");		//(= P2_P1_P1_Flush    0b0)) ;4743
                                        P2_P1_P1_More = 1'b1; $display(";A 4744");		//(= P2_P1_P1_More    0b1)) ;4744
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 4745");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b11101010)) ;4745
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4746");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4746
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4747");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4747
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4748");		//(= P2_P1_P1_Flush    0b0)) ;4748
                                    P2_P1_P1_More = 1'b0; $display(";A 4749");		//(= P2_P1_P1_More    0b0)) ;4749
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 4750");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b10110000)) ;4750
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4751");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4751
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4752");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4752
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4753");		//(= P2_P1_P1_Flush    0b0)) ;4753
                                    P2_P1_P1_More = 1'b0; $display(";A 4754");		//(= P2_P1_P1_More    0b0)) ;4754
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 4755");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b10111000)) ;4755
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 4756");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;4756
                                        P2_P1_P1_EAX <= #1 ((((P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 4758");		//(= P2_P1_P1_EAX    (bv-add (bv-add (bv-add (bv-mul P2_P1_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P1_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P1_P1_InstQueue 0  0b00000000000000000000000100000000)) P2_P1_P1_InstQueue 0 ))) ;4758
                                        P2_P1_P1_More = 1'b0; $display(";A 4759");		//(= P2_P1_P1_More    0b0)) ;4759
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4760");		//(= P2_P1_P1_Flush    0b0)) ;4760
                                        P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 4761");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;4761
                                        P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 4762");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;4762
                                    end
                                    else begin
                                        $display(";A 4757");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;4757
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4763");		//(= P2_P1_P1_Flush    0b0)) ;4763
                                        P2_P1_P1_More = 1'b1; $display(";A 4764");		//(= P2_P1_P1_More    0b1)) ;4764
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 4765");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b10111011)) ;4765
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 4766");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;4766
                                        P2_P1_P1_EBX <= #1 ((((P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P1_P1_InstQueue[((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 4768");		//(= P2_P1_P1_EBX    (bv-add (bv-add (bv-add (bv-mul P2_P1_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P1_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P1_P1_InstQueue 0  0b00000000000000000000000100000000)) P2_P1_P1_InstQueue 0 ))) ;4768
                                        P2_P1_P1_More = 1'b0; $display(";A 4769");		//(= P2_P1_P1_More    0b0)) ;4769
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4770");		//(= P2_P1_P1_Flush    0b0)) ;4770
                                        P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 4771");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;4771
                                        P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 4772");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;4772
                                    end
                                    else begin
                                        $display(";A 4767");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;4767
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4773");		//(= P2_P1_P1_Flush    0b0)) ;4773
                                        P2_P1_P1_More = 1'b1; $display(";A 4774");		//(= P2_P1_P1_More    0b1)) ;4774
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 4775");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b10001011)) ;4775
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 4776");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;4776
                                        if ((P2_P1_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 4778");		//(= (bool-to-bv (bv-slt P2_P1_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;4778
                                            P2_P1_P1_rEIP <= #1 (-P2_P1_P1_EBX); $display(";A 4780");		//(= P2_P1_P1_rEIP    (bv-neg P2_P1_P1_EBX ))) ;4780
                                        end
                                        else begin
                                            $display(";A 4779");		//(= (bool-to-bv (bv-slt P2_P1_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;4779
                                            P2_P1_P1_rEIP <= #1 P2_P1_P1_EBX; $display(";A 4781");		//(= P2_P1_P1_rEIP    P2_P1_P1_EBX )) ;4781
                                        end
                                        P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4782");		//(= P2_P1_P1_RequestPending    0b1)) ;4782
                                        P2_P1_P1_ReadRequest <= #1 1'b1; $display(";A 4783");		//(= P2_P1_P1_ReadRequest    0b1)) ;4783
                                        P2_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 4784");		//(= P2_P1_P1_MemoryFetch    0b1)) ;4784
                                        P2_P1_P1_CodeFetch <= #1 1'b0; $display(";A 4785");		//(= P2_P1_P1_CodeFetch    0b0)) ;4785
                                        if ((P2_P1_P1_READY_n == 1'b0)) begin
                                            $display(";A 4786");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4786
                                            P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4788");		//(= P2_P1_P1_RequestPending    0b0)) ;4788
                                            P2_P1_P1_uWord = (P2_P1_P1_Datai % 32'b00000000000000001000000000000000); $display(";A 4789");		//(= P2_P1_P1_uWord    (bv-smod P2_P1_P1_Datai  0b00000000000000001000000000000000))) ;4789
                                            if ((P2_P1_P1_StateBS16 == 1'b1)) begin
                                                $display(";A 4790");		//(= (bv-comp P2_P1_P1_StateBS16  0b1)   0b1)) ;4790
                                                P2_P1_P1_lWord = (P2_P1_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 4792");		//(= P2_P1_P1_lWord    (bv-smod P2_P1_P1_Datai  0b00000000000000010000000000000000))) ;4792
                                            end
                                            else begin
                                                $display(";A 4791");		//(= (bv-comp P2_P1_P1_StateBS16  0b1)   0b0)) ;4791
                                                P2_P1_P1_rEIP <= #1 (P2_P1_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 4793");		//(= P2_P1_P1_rEIP    (bv-add P2_P1_P1_rEIP  0b00000000000000000000000000000010))) ;4793
                                                P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4794");		//(= P2_P1_P1_RequestPending    0b1)) ;4794
                                                if ((P2_P1_P1_READY_n == 1'b0)) begin
                                                    $display(";A 4795");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4795
                                                    P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4797");		//(= P2_P1_P1_RequestPending    0b0)) ;4797
                                                    P2_P1_P1_lWord = (P2_P1_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 4798");		//(= P2_P1_P1_lWord    (bv-smod P2_P1_P1_Datai  0b00000000000000010000000000000000))) ;4798
                                                end
                                                else begin
                                                    $display(";A 4796");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4796
                                                end
                                            end
                                            if ((P2_P1_P1_READY_n == 1'b0)) begin
                                                $display(";A 4799");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4799
                                                P2_P1_P1_EAX <= #1 ((P2_P1_P1_uWord * 32'b00000000000000010000000000000000) + P2_P1_P1_lWord); $display(";A 4801");		//(= P2_P1_P1_EAX    (bv-add (bv-mul P2_P1_P1_uWord  0b00000000000000010000000000000000) P2_P1_P1_lWord ))) ;4801
                                                P2_P1_P1_More = 1'b0; $display(";A 4802");		//(= P2_P1_P1_More    0b0)) ;4802
                                                P2_P1_P1_Flush = 1'b0; $display(";A 4803");		//(= P2_P1_P1_Flush    0b0)) ;4803
                                                P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4804");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;4804
                                                P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 4805");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;4805
                                            end
                                            else begin
                                                $display(";A 4800");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4800
                                            end
                                        end
                                        else begin
                                            $display(";A 4787");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4787
                                        end
                                    end
                                    else begin
                                        $display(";A 4777");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;4777
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4806");		//(= P2_P1_P1_Flush    0b0)) ;4806
                                        P2_P1_P1_More = 1'b1; $display(";A 4807");		//(= P2_P1_P1_More    0b1)) ;4807
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 4808");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b10001001)) ;4808
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 4809");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;4809
                                        if ((P2_P1_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 4811");		//(= (bool-to-bv (bv-slt P2_P1_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;4811
                                            P2_P1_P1_rEIP <= #1 P2_P1_P1_EBX; $display(";A 4813");		//(= P2_P1_P1_rEIP    P2_P1_P1_EBX )) ;4813
                                        end
                                        else begin
                                            $display(";A 4812");		//(= (bool-to-bv (bv-slt P2_P1_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;4812
                                            P2_P1_P1_rEIP <= #1 P2_P1_P1_EBX; $display(";A 4814");		//(= P2_P1_P1_rEIP    P2_P1_P1_EBX )) ;4814
                                        end
                                        P2_P1_P1_lWord = (P2_P1_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 4815");		//(= P2_P1_P1_lWord    (bv-smod P2_P1_P1_EAX  0b00000000000000010000000000000000))) ;4815
                                        P2_P1_P1_uWord = ((P2_P1_P1_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 4816");		//(= P2_P1_P1_uWord    (bv-smod (bv-sdiv P2_P1_P1_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;4816
                                        P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4817");		//(= P2_P1_P1_RequestPending    0b1)) ;4817
                                        P2_P1_P1_ReadRequest <= #1 1'b0; $display(";A 4818");		//(= P2_P1_P1_ReadRequest    0b0)) ;4818
                                        P2_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 4819");		//(= P2_P1_P1_MemoryFetch    0b1)) ;4819
                                        P2_P1_P1_CodeFetch <= #1 1'b0; $display(";A 4820");		//(= P2_P1_P1_CodeFetch    0b0)) ;4820
                                        if (((P2_P1_P1_State == 32'b00000000000000000000000000000010) | (P2_P1_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 4821");		//(= (bv-or (bv-comp P2_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P1_State  0b00000000000000000000000000000100))   0b1)) ;4821
                                            P2_P1_P1_Datao <= #1 ((P2_P1_P1_uWord * 32'b00000000000000010000000000000000) + P2_P1_P1_lWord); $display(";A 4823");		//(= P2_P1_P1_Datao    (bv-add (bv-mul P2_P1_P1_uWord  0b00000000000000010000000000000000) P2_P1_P1_lWord ))) ;4823
                                            if ((P2_P1_P1_READY_n == 1'b0)) begin
                                                $display(";A 4824");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4824
                                                P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4826");		//(= P2_P1_P1_RequestPending    0b0)) ;4826
                                                if ((P2_P1_P1_StateBS16 == 1'b0)) begin
                                                    $display(";A 4827");		//(= (bv-comp P2_P1_P1_StateBS16  0b0)   0b1)) ;4827
                                                    P2_P1_P1_rEIP <= #1 (P2_P1_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 4829");		//(= P2_P1_P1_rEIP    (bv-add P2_P1_P1_rEIP  0b00000000000000000000000000000010))) ;4829
                                                    P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4830");		//(= P2_P1_P1_RequestPending    0b1)) ;4830
                                                    P2_P1_P1_ReadRequest <= #1 1'b0; $display(";A 4831");		//(= P2_P1_P1_ReadRequest    0b0)) ;4831
                                                    P2_P1_P1_MemoryFetch <= #1 1'b1; $display(";A 4832");		//(= P2_P1_P1_MemoryFetch    0b1)) ;4832
                                                    P2_P1_P1_CodeFetch <= #1 1'b0; $display(";A 4833");		//(= P2_P1_P1_CodeFetch    0b0)) ;4833
                                                    P2_P1_P1_State2 = 4'sb0110; $display(";A 4834");		//(= P2_P1_P1_State2    0b0110)) ;4834
                                                end
                                                else begin
                                                    $display(";A 4828");		//(= (bv-comp P2_P1_P1_StateBS16  0b0)   0b0)) ;4828
                                                end
                                                P2_P1_P1_More = 1'b0; $display(";A 4835");		//(= P2_P1_P1_More    0b0)) ;4835
                                                P2_P1_P1_Flush = 1'b0; $display(";A 4836");		//(= P2_P1_P1_Flush    0b0)) ;4836
                                                P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4837");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;4837
                                                P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 4838");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;4838
                                            end
                                            else begin
                                                $display(";A 4825");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4825
                                            end
                                        end
                                        else begin
                                            $display(";A 4822");		//(= (bv-or (bv-comp P2_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P1_State  0b00000000000000000000000000000100))   0b0)) ;4822
                                        end
                                    end
                                    else begin
                                        $display(";A 4810");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;4810
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4839");		//(= P2_P1_P1_Flush    0b0)) ;4839
                                        P2_P1_P1_More = 1'b1; $display(";A 4840");		//(= P2_P1_P1_More    0b1)) ;4840
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 4841");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b11100100)) ;4841
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 4842");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;4842
                                        P2_P1_P1_rEIP <= #1 (P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 4844");		//(= P2_P1_P1_rEIP    (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;4844
                                        P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4845");		//(= P2_P1_P1_RequestPending    0b1)) ;4845
                                        P2_P1_P1_ReadRequest <= #1 1'b1; $display(";A 4846");		//(= P2_P1_P1_ReadRequest    0b1)) ;4846
                                        P2_P1_P1_MemoryFetch <= #1 1'b0; $display(";A 4847");		//(= P2_P1_P1_MemoryFetch    0b0)) ;4847
                                        P2_P1_P1_CodeFetch <= #1 1'b0; $display(";A 4848");		//(= P2_P1_P1_CodeFetch    0b0)) ;4848
                                        if ((P2_P1_P1_READY_n == 1'b0)) begin
                                            $display(";A 4849");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4849
                                            P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4851");		//(= P2_P1_P1_RequestPending    0b0)) ;4851
                                            P2_P1_P1_EAX <= #1 P2_P1_P1_Datai; $display(";A 4852");		//(= P2_P1_P1_EAX    P2_P1_P1_Datai )) ;4852
                                            P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4853");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;4853
                                            P2_P1_P1_InstQueueRd_Addr = (P2_P1_P1_InstQueueRd_Addr + 5'b00010); $display(";A 4854");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-add P2_P1_P1_InstQueueRd_Addr  0b00010))) ;4854
                                            P2_P1_P1_Flush = 1'b0; $display(";A 4855");		//(= P2_P1_P1_Flush    0b0)) ;4855
                                            P2_P1_P1_More = 1'b0; $display(";A 4856");		//(= P2_P1_P1_More    0b0)) ;4856
                                        end
                                        else begin
                                            $display(";A 4850");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4850
                                        end
                                    end
                                    else begin
                                        $display(";A 4843");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;4843
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4857");		//(= P2_P1_P1_Flush    0b0)) ;4857
                                        P2_P1_P1_More = 1'b1; $display(";A 4858");		//(= P2_P1_P1_More    0b1)) ;4858
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 4859");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b11100110)) ;4859
                                    if (((P2_P1_P1_InstQueueWr_Addr - P2_P1_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 4860");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;4860
                                        P2_P1_P1_rEIP <= #1 (P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 4862");		//(= P2_P1_P1_rEIP    (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;4862
                                        P2_P1_P1_RequestPending <= #1 1'b1; $display(";A 4863");		//(= P2_P1_P1_RequestPending    0b1)) ;4863
                                        P2_P1_P1_ReadRequest <= #1 1'b0; $display(";A 4864");		//(= P2_P1_P1_ReadRequest    0b0)) ;4864
                                        P2_P1_P1_MemoryFetch <= #1 1'b0; $display(";A 4865");		//(= P2_P1_P1_MemoryFetch    0b0)) ;4865
                                        P2_P1_P1_CodeFetch <= #1 1'b0; $display(";A 4866");		//(= P2_P1_P1_CodeFetch    0b0)) ;4866
                                        if (((P2_P1_P1_State == 32'b00000000000000000000000000000010) | (P2_P1_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 4867");		//(= (bv-or (bv-comp P2_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P1_State  0b00000000000000000000000000000100))   0b1)) ;4867
                                            P2_P1_P1_fWord = (P2_P1_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 4869");		//(= P2_P1_P1_fWord    (bv-smod P2_P1_P1_EAX  0b00000000000000010000000000000000))) ;4869
                                            P2_P1_P1_Datao <= #1 P2_P1_P1_fWord; $display(";A 4870");		//(= P2_P1_P1_Datao    P2_P1_P1_fWord )) ;4870
                                            if ((P2_P1_P1_READY_n == 1'b0)) begin
                                                $display(";A 4871");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4871
                                                P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4873");		//(= P2_P1_P1_RequestPending    0b0)) ;4873
                                                P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4874");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;4874
                                                P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 4875");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;4875
                                                P2_P1_P1_Flush = 1'b0; $display(";A 4876");		//(= P2_P1_P1_Flush    0b0)) ;4876
                                                P2_P1_P1_More = 1'b0; $display(";A 4877");		//(= P2_P1_P1_More    0b0)) ;4877
                                            end
                                            else begin
                                                $display(";A 4872");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4872
                                            end
                                        end
                                        else begin
                                            $display(";A 4868");		//(= (bv-or (bv-comp P2_P1_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P1_State  0b00000000000000000000000000000100))   0b0)) ;4868
                                        end
                                    end
                                    else begin
                                        $display(";A 4861");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P1_InstQueueWr_Addr  P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;4861
                                        P2_P1_P1_Flush = 1'b0; $display(";A 4878");		//(= P2_P1_P1_Flush    0b0)) ;4878
                                        P2_P1_P1_More = 1'b1; $display(";A 4879");		//(= P2_P1_P1_More    0b1)) ;4879
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 4880");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b00000100)) ;4880
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4881");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4881
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4882");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4882
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4883");		//(= P2_P1_P1_Flush    0b0)) ;4883
                                    P2_P1_P1_More = 1'b0; $display(";A 4884");		//(= P2_P1_P1_More    0b0)) ;4884
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 4885");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b00000101)) ;4885
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4886");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4886
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4887");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4887
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4888");		//(= P2_P1_P1_Flush    0b0)) ;4888
                                    P2_P1_P1_More = 1'b0; $display(";A 4889");		//(= P2_P1_P1_More    0b0)) ;4889
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 4890");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b11010000)) ;4890
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4891");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;4891
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 4892");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;4892
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4893");		//(= P2_P1_P1_Flush    0b0)) ;4893
                                    P2_P1_P1_More = 1'b0; $display(";A 4894");		//(= P2_P1_P1_More    0b0)) ;4894
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 4895");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b11000000)) ;4895
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 4896");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;4896
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 4897");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;4897
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4898");		//(= P2_P1_P1_Flush    0b0)) ;4898
                                    P2_P1_P1_More = 1'b0; $display(";A 4899");		//(= P2_P1_P1_More    0b0)) ;4899
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 4900");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b01000000)) ;4900
                                    P2_P1_P1_EAX <= #1 (P2_P1_P1_EAX + 32'sb00000000000000000000000000000001); $display(";A 4901");		//(= P2_P1_P1_EAX    (bv-add P2_P1_P1_EAX  0b00000000000000000000000000000001))) ;4901
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4902");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4902
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4903");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4903
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4904");		//(= P2_P1_P1_Flush    0b0)) ;4904
                                    P2_P1_P1_More = 1'b0; $display(";A 4905");		//(= P2_P1_P1_More    0b0)) ;4905
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 4906");		//(= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr )   0b01000011)) ;4906
                                    P2_P1_P1_EBX <= #1 (P2_P1_P1_EBX + 32'sb00000000000000000000000000000001); $display(";A 4907");		//(= P2_P1_P1_EBX    (bv-add P2_P1_P1_EBX  0b00000000000000000000000000000001))) ;4907
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4908");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4908
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4909");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4909
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4910");		//(= P2_P1_P1_Flush    0b0)) ;4910
                                    P2_P1_P1_More = 1'b0; $display(";A 4911");		//(= P2_P1_P1_More    0b0)) ;4911
                                end
                            default:
                                begin
                                    $display(";A 4912");		//(= (and (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b10010000) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b01100110) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b11101011) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b11101001) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b11101010) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b10110000) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b10111000) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b10111011) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b10001011) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b10001001) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b11100100) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b11100110) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b00000100) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b00000101) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b11010000) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b11000000) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b01000000) (/= ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ) 0b01000011))   true)) ;4912
                                    P2_P1_P1_InstAddrPointer = (P2_P1_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 4913");		//(= P2_P1_P1_InstAddrPointer    (bv-add P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;4913
                                    P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4914");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4914
                                    P2_P1_P1_Flush = 1'b0; $display(";A 4915");		//(= P2_P1_P1_Flush    0b0)) ;4915
                                    P2_P1_P1_More = 1'b0; $display(";A 4916");		//(= P2_P1_P1_More    0b0)) ;4916
                                end
                        endcase
                        if (((~(P2_P1_P1_InstQueueRd_Addr < P2_P1_P1_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P2_P1_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P2_P1_P1_Flush) | P2_P1_P1_More))) begin
                            $display(";A 4917");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P1_P1_InstQueueRd_Addr  P2_P1_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P1_P1_Flush ) P2_P1_P1_More ))   0b1)) ;4917
                            P2_P1_P1_State2 = 4'sb0111; $display(";A 4919");		//(= P2_P1_P1_State2    0b0111)) ;4919
                        end
                        else begin
                            $display(";A 4918");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P1_P1_InstQueueRd_Addr  P2_P1_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P1_P1_Flush ) P2_P1_P1_More ))   0b0)) ;4918
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 4920");		//(= P2_P1_P1_State2    0b0110)) ;4920
                        P2_P1_P1_Datao <= #1 ((P2_P1_P1_uWord * 32'b00000000000000010000000000000000) + P2_P1_P1_lWord); $display(";A 4921");		//(= P2_P1_P1_Datao    (bv-add (bv-mul P2_P1_P1_uWord  0b00000000000000010000000000000000) P2_P1_P1_lWord ))) ;4921
                        if ((P2_P1_P1_READY_n == 1'b0)) begin
                            $display(";A 4922");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b1)) ;4922
                            P2_P1_P1_RequestPending <= #1 1'b0; $display(";A 4924");		//(= P2_P1_P1_RequestPending    0b0)) ;4924
                            P2_P1_P1_State2 = 4'sb0101; $display(";A 4925");		//(= P2_P1_P1_State2    0b0101)) ;4925
                        end
                        else begin
                            $display(";A 4923");		//(= (bv-comp P2_P1_P1_READY_n  0b0)   0b0)) ;4923
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 4926");		//(= P2_P1_P1_State2    0b0111)) ;4926
                        if (P2_P1_P1_Flush) begin
                            $display(";A 4927");		//(= P2_P1_P1_Flush    0b1)) ;4927
                            P2_P1_P1_InstQueueRd_Addr = 5'sb00001; $display(";A 4929");		//(= P2_P1_P1_InstQueueRd_Addr    0b00001)) ;4929
                            P2_P1_P1_InstQueueWr_Addr = 5'sb00001; $display(";A 4930");		//(= P2_P1_P1_InstQueueWr_Addr    0b00001)) ;4930
                            if ((P2_P1_P1_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 4931");		//(= (bool-to-bv (bv-slt P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;4931
                                P2_P1_P1_fWord = (-P2_P1_P1_InstAddrPointer); $display(";A 4933");		//(= P2_P1_P1_fWord    (bv-neg P2_P1_P1_InstAddrPointer ))) ;4933
                            end
                            else begin
                                $display(";A 4932");		//(= (bool-to-bv (bv-slt P2_P1_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;4932
                                P2_P1_P1_fWord = P2_P1_P1_InstAddrPointer; $display(";A 4934");		//(= P2_P1_P1_fWord    P2_P1_P1_InstAddrPointer )) ;4934
                            end
                            if (((P2_P1_P1_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 4935");		//(= (bv-comp (bv-smod P2_P1_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;4935
                                P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + (P2_P1_P1_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 4937");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  (bv-smod P2_P1_P1_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;4937
                            end
                            else begin
                                $display(";A 4936");		//(= (bv-comp (bv-smod P2_P1_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;4936
                            end
                        end
                        else begin
                            $display(";A 4928");		//(= P2_P1_P1_Flush    0b0)) ;4928
                        end
                        if (((32'b00000000000000000000000000001111 - P2_P1_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 4938");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;4938
                            P2_P1_P1_State2 = 4'sb1000; $display(";A 4940");		//(= P2_P1_P1_State2    0b1000)) ;4940
                            P2_P1_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 4941");		//(= P2_P1_P1_InstQueueWr_Addr    0b00000)) ;4941
                        end
                        else begin
                            $display(";A 4939");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;4939
                            P2_P1_P1_State2 = 4'sb1001; $display(";A 4942");		//(= P2_P1_P1_State2    0b1001)) ;4942
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 4943");		//(= P2_P1_P1_State2    0b1000)) ;4943
                        if ((P2_P1_P1_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 4944");		//(= (bool-to-bv (bv-le P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;4944
                            P2_P1_P1_InstQueue[P2_P1_P1_InstQueueWr_Addr] = P2_P1_P1_InstQueue[P2_P1_P1_InstQueueRd_Addr]; $display(";A 4946");		//(= P2_P1_P1_InstQueue    ( P2_P1_P1_InstQueue P2_P1_P1_InstQueueRd_Addr ))) ;4946
                            P2_P1_P1_InstQueueRd_Addr = ((P2_P1_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4947");		//(= P2_P1_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4947
                            P2_P1_P1_InstQueueWr_Addr = ((P2_P1_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 4948");		//(= P2_P1_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;4948
                            P2_P1_P1_State2 = 4'sb1000; $display(";A 4949");		//(= P2_P1_P1_State2    0b1000)) ;4949
                        end
                        else begin
                            $display(";A 4945");		//(= (bool-to-bv (bv-le P2_P1_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;4945
                            P2_P1_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 4950");		//(= P2_P1_P1_InstQueueRd_Addr    0b00000)) ;4950
                            P2_P1_P1_State2 = 4'sb1001; $display(";A 4951");		//(= P2_P1_P1_State2    0b1001)) ;4951
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 4952");		//(= P2_P1_P1_State2    0b1001)) ;4952
                        P2_P1_P1_rEIP <= #1 P2_P1_P1_PhyAddrPointer; $display(";A 4953");		//(= P2_P1_P1_rEIP    P2_P1_P1_PhyAddrPointer )) ;4953
                        P2_P1_P1_State2 = 4'sb0001; $display(";A 4954");		//(= P2_P1_P1_State2    0b0001)) ;4954
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:7474
    always @(posedge P2_P1_P1_RESET or posedge P2_P1_P1_CLOCK) begin
        if ((P2_P1_P1_RESET == 1'b1)) begin
            $display(";A 4955");		//(= (bv-comp P2_P1_P1_RESET  0b1)   0b1)) ;4955
            P2_P1_P1_ByteEnable <= #1 4'b0000; $display(";A 4957");		//(= P2_P1_P1_ByteEnable    0b0000)) ;4957
            P2_P1_P1_NonAligned <= #1 1'b0; $display(";A 4958");		//(= P2_P1_P1_NonAligned    0b0)) ;4958
        end
        else begin
            $display(";A 4956");		//(= (bv-comp P2_P1_P1_RESET  0b1)   0b0)) ;4956
            case (P2_P1_P1_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 4959");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000000)) ;4959
                        case ((P2_P1_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 4960");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;4960
                                    P2_P1_P1_ByteEnable <= #1 4'b1110; $display(";A 4961");		//(= P2_P1_P1_ByteEnable    0b1110)) ;4961
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 4962");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;4962
                                    P2_P1_P1_ByteEnable <= #1 4'b1101; $display(";A 4963");		//(= P2_P1_P1_ByteEnable    0b1101)) ;4963
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 4964");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;4964
                                    P2_P1_P1_ByteEnable <= #1 4'b1011; $display(";A 4965");		//(= P2_P1_P1_ByteEnable    0b1011)) ;4965
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 4966");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;4966
                                    P2_P1_P1_ByteEnable <= #1 4'b0111; $display(";A 4967");		//(= P2_P1_P1_ByteEnable    0b0111)) ;4967
                                end
                            default:
                                begin
                                    $display(";A 4968");		//(= (and (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;4968
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 4969");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000001)) ;4969
                        case ((P2_P1_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 4970");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;4970
                                    P2_P1_P1_ByteEnable <= #1 4'b1100; $display(";A 4971");		//(= P2_P1_P1_ByteEnable    0b1100)) ;4971
                                    P2_P1_P1_NonAligned <= #1 1'b0; $display(";A 4972");		//(= P2_P1_P1_NonAligned    0b0)) ;4972
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 4973");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;4973
                                    P2_P1_P1_ByteEnable <= #1 4'b1001; $display(";A 4974");		//(= P2_P1_P1_ByteEnable    0b1001)) ;4974
                                    P2_P1_P1_NonAligned <= #1 1'b0; $display(";A 4975");		//(= P2_P1_P1_NonAligned    0b0)) ;4975
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 4976");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;4976
                                    P2_P1_P1_ByteEnable <= #1 4'b0011; $display(";A 4977");		//(= P2_P1_P1_ByteEnable    0b0011)) ;4977
                                    P2_P1_P1_NonAligned <= #1 1'b0; $display(";A 4978");		//(= P2_P1_P1_NonAligned    0b0)) ;4978
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 4979");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;4979
                                    P2_P1_P1_ByteEnable <= #1 4'b0111; $display(";A 4980");		//(= P2_P1_P1_ByteEnable    0b0111)) ;4980
                                    P2_P1_P1_NonAligned <= #1 1'b1; $display(";A 4981");		//(= P2_P1_P1_NonAligned    0b1)) ;4981
                                end
                            default:
                                begin
                                    $display(";A 4982");		//(= (and (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;4982
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 4983");		//(= P2_P1_P1_DataWidth    0b00000000000000000000000000000010)) ;4983
                        case ((P2_P1_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 4984");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;4984
                                    P2_P1_P1_ByteEnable <= #1 4'b0000; $display(";A 4985");		//(= P2_P1_P1_ByteEnable    0b0000)) ;4985
                                    P2_P1_P1_NonAligned <= #1 1'b0; $display(";A 4986");		//(= P2_P1_P1_NonAligned    0b0)) ;4986
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 4987");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;4987
                                    P2_P1_P1_ByteEnable <= #1 4'b0001; $display(";A 4988");		//(= P2_P1_P1_ByteEnable    0b0001)) ;4988
                                    P2_P1_P1_NonAligned <= #1 1'b1; $display(";A 4989");		//(= P2_P1_P1_NonAligned    0b1)) ;4989
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 4990");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;4990
                                    P2_P1_P1_NonAligned <= #1 1'b1; $display(";A 4991");		//(= P2_P1_P1_NonAligned    0b1)) ;4991
                                    P2_P1_P1_ByteEnable <= #1 4'b0011; $display(";A 4992");		//(= P2_P1_P1_ByteEnable    0b0011)) ;4992
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 4993");		//(= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;4993
                                    P2_P1_P1_NonAligned <= #1 1'b1; $display(";A 4994");		//(= P2_P1_P1_NonAligned    0b1)) ;4994
                                    P2_P1_P1_ByteEnable <= #1 4'b0111; $display(";A 4995");		//(= P2_P1_P1_ByteEnable    0b0111)) ;4995
                                end
                            default:
                                begin
                                    $display(";A 4996");		//(= (and (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;4996
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 4997");		//(= (and (/= P2_P1_P1_DataWidth  0b00000000000000000000000000000000) (/= P2_P1_P1_DataWidth  0b00000000000000000000000000000001) (/= P2_P1_P1_DataWidth  0b00000000000000000000000000000010))   true)) ;4997
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:7662
    always @(posedge P2_P1_P2_RESET or posedge P2_P1_P2_CLOCK) begin
        if ((P2_P1_P2_RESET == 1'b1)) begin
            $display(";A 4998");		//(= (bv-comp P2_P1_P2_RESET  0b1)   0b1)) ;4998
            P2_P1_P2_BE_n <= #1 4'b0000; $display(";A 5000");		//(= P2_P1_P2_BE_n    0b0000)) ;5000
            P2_P1_P2_Address <= #1 30'sb000000000000000000000000000000; $display(";A 5001");		//(= P2_P1_P2_Address    0b000000000000000000000000000000)) ;5001
            P2_P1_P2_W_R_n <= #1 1'b0; $display(";A 5002");		//(= P2_P1_P2_W_R_n    0b0)) ;5002
            P2_P1_P2_D_C_n <= #1 1'b0; $display(";A 5003");		//(= P2_P1_P2_D_C_n    0b0)) ;5003
            P2_P1_P2_M_IO_n <= #1 1'b0; $display(";A 5004");		//(= P2_P1_P2_M_IO_n    0b0)) ;5004
            P2_P1_P2_ADS_n <= #1 1'b0; $display(";A 5005");		//(= P2_P1_P2_ADS_n    0b0)) ;5005
            P2_P1_P2_State <= #1 3'sb000; $display(";A 5006");		//(= P2_P1_P2_State    0b000)) ;5006
            P2_P1_P2_StateNA <= #1 1'b0; $display(";A 5007");		//(= P2_P1_P2_StateNA    0b0)) ;5007
            P2_P1_P2_StateBS16 <= #1 1'b0; $display(";A 5008");		//(= P2_P1_P2_StateBS16    0b0)) ;5008
            P2_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 5009");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000000)) ;5009
        end
        else begin
            $display(";A 4999");		//(= (bv-comp P2_P1_P2_RESET  0b1)   0b0)) ;4999
            case (P2_P1_P2_State)
                3'b000 :
                    begin
                        $display(";A 5010");		//(= P2_P1_P2_State    0b000)) ;5010
                        P2_P1_P2_D_C_n <= #1 1'b1; $display(";A 5011");		//(= P2_P1_P2_D_C_n    0b1)) ;5011
                        P2_P1_P2_ADS_n <= #1 1'b1; $display(";A 5012");		//(= P2_P1_P2_ADS_n    0b1)) ;5012
                        P2_P1_P2_State <= #1 3'sb001; $display(";A 5013");		//(= P2_P1_P2_State    0b001)) ;5013
                        P2_P1_P2_StateNA <= #1 1'b1; $display(";A 5014");		//(= P2_P1_P2_StateNA    0b1)) ;5014
                        P2_P1_P2_StateBS16 <= #1 1'b1; $display(";A 5015");		//(= P2_P1_P2_StateBS16    0b1)) ;5015
                        P2_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 5016");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;5016
                        P2_P1_P2_State <= #1 3'sb001; $display(";A 5017");		//(= P2_P1_P2_State    0b001)) ;5017
                    end
                3'b001 :
                    begin
                        $display(";A 5018");		//(= P2_P1_P2_State    0b001)) ;5018
                        if ((P2_P1_P2_RequestPending == 1'b1)) begin
                            $display(";A 5019");		//(= (bv-comp P2_P1_P2_RequestPending  0b1)   0b1)) ;5019
                            P2_P1_P2_State <= #1 3'sb010; $display(";A 5021");		//(= P2_P1_P2_State    0b010)) ;5021
                        end
                        else begin
                            $display(";A 5020");		//(= (bv-comp P2_P1_P2_RequestPending  0b1)   0b0)) ;5020
                            if ((P2_P1_P2_HOLD == 1'b1)) begin
                                $display(";A 5022");		//(= (bv-comp P2_P1_P2_HOLD  0b1)   0b1)) ;5022
                                P2_P1_P2_State <= #1 3'sb101; $display(";A 5024");		//(= P2_P1_P2_State    0b101)) ;5024
                            end
                            else begin
                                $display(";A 5023");		//(= (bv-comp P2_P1_P2_HOLD  0b1)   0b0)) ;5023
                                P2_P1_P2_State <= #1 3'sb001; $display(";A 5025");		//(= P2_P1_P2_State    0b001)) ;5025
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 5026");		//(= P2_P1_P2_State    0b010)) ;5026
                        P2_P1_P2_Address <= #1 ((P2_P1_P2_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 5027");		//(= P2_P1_P2_Address    (bv-smod (bv-sdiv P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;5027
                        P2_P1_P2_BE_n <= #1 P2_P1_P2_ByteEnable; $display(";A 5028");		//(= P2_P1_P2_BE_n    P2_P1_P2_ByteEnable )) ;5028
                        P2_P1_P2_M_IO_n <= #1 P2_P1_P2_MemoryFetch; $display(";A 5029");		//(= P2_P1_P2_M_IO_n    P2_P1_P2_MemoryFetch )) ;5029
                        if ((P2_P1_P2_ReadRequest == 1'b1)) begin
                            $display(";A 5030");		//(= (bv-comp P2_P1_P2_ReadRequest  0b1)   0b1)) ;5030
                            P2_P1_P2_W_R_n <= #1 1'b0; $display(";A 5032");		//(= P2_P1_P2_W_R_n    0b0)) ;5032
                        end
                        else begin
                            $display(";A 5031");		//(= (bv-comp P2_P1_P2_ReadRequest  0b1)   0b0)) ;5031
                            P2_P1_P2_W_R_n <= #1 1'b1; $display(";A 5033");		//(= P2_P1_P2_W_R_n    0b1)) ;5033
                        end
                        if ((P2_P1_P2_CodeFetch == 1'b1)) begin
                            $display(";A 5034");		//(= (bv-comp P2_P1_P2_CodeFetch  0b1)   0b1)) ;5034
                            P2_P1_P2_D_C_n <= #1 1'b0; $display(";A 5036");		//(= P2_P1_P2_D_C_n    0b0)) ;5036
                        end
                        else begin
                            $display(";A 5035");		//(= (bv-comp P2_P1_P2_CodeFetch  0b1)   0b0)) ;5035
                            P2_P1_P2_D_C_n <= #1 1'b1; $display(";A 5037");		//(= P2_P1_P2_D_C_n    0b1)) ;5037
                        end
                        P2_P1_P2_ADS_n <= #1 1'b0; $display(";A 5038");		//(= P2_P1_P2_ADS_n    0b0)) ;5038
                        P2_P1_P2_State <= #1 3'sb011; $display(";A 5039");		//(= P2_P1_P2_State    0b011)) ;5039
                    end
                3'b011 :
                    begin
                        $display(";A 5040");		//(= P2_P1_P2_State    0b011)) ;5040
                        if ((((P2_P1_P2_READY_n == 1'b0) & (P2_P1_P2_HOLD == 1'b0)) & (P2_P1_P2_RequestPending == 1'b1))) begin
                            $display(";A 5041");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b1))   0b1)) ;5041
                            P2_P1_P2_State <= #1 3'sb010; $display(";A 5043");		//(= P2_P1_P2_State    0b010)) ;5043
                        end
                        else begin
                            $display(";A 5042");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b1))   0b0)) ;5042
                            if (((P2_P1_P2_READY_n == 1'b1) & (P2_P1_P2_NA_n == 1'b1))) begin
                                $display(";A 5044");		//(= (bv-and (bv-comp P2_P1_P2_READY_n  0b1) (bv-comp P2_P1_P2_NA_n  0b1))   0b1)) ;5044
                            end
                            else begin
                                $display(";A 5045");		//(= (bv-and (bv-comp P2_P1_P2_READY_n  0b1) (bv-comp P2_P1_P2_NA_n  0b1))   0b0)) ;5045
                                if ((((P2_P1_P2_RequestPending == 1'b1) | (P2_P1_P2_HOLD == 1'b1)) & ((P2_P1_P2_READY_n == 1'b1) & (P2_P1_P2_NA_n == 1'b0)))) begin
                                    $display(";A 5046");		//(= (bv-and (bv-or (bv-comp P2_P1_P2_RequestPending  0b1) (bv-comp P2_P1_P2_HOLD  0b1)) (bv-and (bv-comp P2_P1_P2_READY_n  0b1) (bv-comp P2_P1_P2_NA_n  0b0)))   0b1)) ;5046
                                    P2_P1_P2_State <= #1 3'sb111; $display(";A 5048");		//(= P2_P1_P2_State    0b111)) ;5048
                                end
                                else begin
                                    $display(";A 5047");		//(= (bv-and (bv-or (bv-comp P2_P1_P2_RequestPending  0b1) (bv-comp P2_P1_P2_HOLD  0b1)) (bv-and (bv-comp P2_P1_P2_READY_n  0b1) (bv-comp P2_P1_P2_NA_n  0b0)))   0b0)) ;5047
                                    if (((((P2_P1_P2_RequestPending == 1'b1) & (P2_P1_P2_HOLD == 1'b0)) & (P2_P1_P2_READY_n == 1'b1)) & (P2_P1_P2_NA_n == 1'b0))) begin
                                        $display(";A 5049");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P1_P2_RequestPending  0b1) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_READY_n  0b1)) (bv-comp P2_P1_P2_NA_n  0b0))   0b1)) ;5049
                                        P2_P1_P2_State <= #1 3'sb110; $display(";A 5051");		//(= P2_P1_P2_State    0b110)) ;5051
                                    end
                                    else begin
                                        $display(";A 5050");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P1_P2_RequestPending  0b1) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_READY_n  0b1)) (bv-comp P2_P1_P2_NA_n  0b0))   0b0)) ;5050
                                        if ((((P2_P1_P2_RequestPending == 1'b0) & (P2_P1_P2_HOLD == 1'b0)) & (P2_P1_P2_READY_n == 1'b0))) begin
                                            $display(";A 5052");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_RequestPending  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_READY_n  0b0))   0b1)) ;5052
                                            P2_P1_P2_State <= #1 3'sb001; $display(";A 5054");		//(= P2_P1_P2_State    0b001)) ;5054
                                        end
                                        else begin
                                            $display(";A 5053");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_RequestPending  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_READY_n  0b0))   0b0)) ;5053
                                            if (((P2_P1_P2_HOLD == 1'b1) & (P2_P1_P2_READY_n == 1'b1))) begin
                                                $display(";A 5055");		//(= (bv-and (bv-comp P2_P1_P2_HOLD  0b1) (bv-comp P2_P1_P2_READY_n  0b1))   0b1)) ;5055
                                                P2_P1_P2_State <= #1 3'sb101; $display(";A 5057");		//(= P2_P1_P2_State    0b101)) ;5057
                                            end
                                            else begin
                                                $display(";A 5056");		//(= (bv-and (bv-comp P2_P1_P2_HOLD  0b1) (bv-comp P2_P1_P2_READY_n  0b1))   0b0)) ;5056
                                                P2_P1_P2_State <= #1 3'sb011; $display(";A 5058");		//(= P2_P1_P2_State    0b011)) ;5058
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P2_P1_P2_StateBS16 <= #1 P2_P1_P2_BS16_n; $display(";A 5059");		//(= P2_P1_P2_StateBS16    P2_P1_P2_BS16_n )) ;5059
                        if ((P2_P1_P2_BS16_n == 1'b0)) begin
                            $display(";A 5060");		//(= (bv-comp P2_P1_P2_BS16_n  0b0)   0b1)) ;5060
                            P2_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 5062");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000001)) ;5062
                        end
                        else begin
                            $display(";A 5061");		//(= (bv-comp P2_P1_P2_BS16_n  0b0)   0b0)) ;5061
                            P2_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 5063");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;5063
                        end
                        P2_P1_P2_StateNA <= #1 P2_P1_P2_NA_n; $display(";A 5064");		//(= P2_P1_P2_StateNA    P2_P1_P2_NA_n )) ;5064
                        P2_P1_P2_ADS_n <= #1 1'b1; $display(";A 5065");		//(= P2_P1_P2_ADS_n    0b1)) ;5065
                    end
                3'b100 :
                    begin
                        $display(";A 5066");		//(= P2_P1_P2_State    0b100)) ;5066
                        if ((((P2_P1_P2_NA_n == 1'b0) & (P2_P1_P2_HOLD == 1'b0)) & (P2_P1_P2_RequestPending == 1'b1))) begin
                            $display(";A 5067");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_NA_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b1))   0b1)) ;5067
                            P2_P1_P2_State <= #1 3'sb110; $display(";A 5069");		//(= P2_P1_P2_State    0b110)) ;5069
                        end
                        else begin
                            $display(";A 5068");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_NA_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b1))   0b0)) ;5068
                            if (((P2_P1_P2_NA_n == 1'b0) & ((P2_P1_P2_HOLD == 1'b1) | (P2_P1_P2_RequestPending == 1'b0)))) begin
                                $display(";A 5070");		//(= (bv-and (bv-comp P2_P1_P2_NA_n  0b0) (bv-or (bv-comp P2_P1_P2_HOLD  0b1) (bv-comp P2_P1_P2_RequestPending  0b0)))   0b1)) ;5070
                                P2_P1_P2_State <= #1 3'sb111; $display(";A 5072");		//(= P2_P1_P2_State    0b111)) ;5072
                            end
                            else begin
                                $display(";A 5071");		//(= (bv-and (bv-comp P2_P1_P2_NA_n  0b0) (bv-or (bv-comp P2_P1_P2_HOLD  0b1) (bv-comp P2_P1_P2_RequestPending  0b0)))   0b0)) ;5071
                                if ((P2_P1_P2_NA_n == 1'b1)) begin
                                    $display(";A 5073");		//(= (bv-comp P2_P1_P2_NA_n  0b1)   0b1)) ;5073
                                    P2_P1_P2_State <= #1 3'sb011; $display(";A 5075");		//(= P2_P1_P2_State    0b011)) ;5075
                                end
                                else begin
                                    $display(";A 5074");		//(= (bv-comp P2_P1_P2_NA_n  0b1)   0b0)) ;5074
                                    P2_P1_P2_State <= #1 3'sb100; $display(";A 5076");		//(= P2_P1_P2_State    0b100)) ;5076
                                end
                            end
                        end
                        P2_P1_P2_StateBS16 <= #1 P2_P1_P2_BS16_n; $display(";A 5077");		//(= P2_P1_P2_StateBS16    P2_P1_P2_BS16_n )) ;5077
                        if ((P2_P1_P2_BS16_n == 1'b0)) begin
                            $display(";A 5078");		//(= (bv-comp P2_P1_P2_BS16_n  0b0)   0b1)) ;5078
                            P2_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 5080");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000001)) ;5080
                        end
                        else begin
                            $display(";A 5079");		//(= (bv-comp P2_P1_P2_BS16_n  0b0)   0b0)) ;5079
                            P2_P1_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 5081");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;5081
                        end
                        P2_P1_P2_StateNA <= #1 P2_P1_P2_NA_n; $display(";A 5082");		//(= P2_P1_P2_StateNA    P2_P1_P2_NA_n )) ;5082
                        P2_P1_P2_ADS_n <= #1 1'b1; $display(";A 5083");		//(= P2_P1_P2_ADS_n    0b1)) ;5083
                    end
                3'b101 :
                    begin
                        $display(";A 5084");		//(= P2_P1_P2_State    0b101)) ;5084
                        if (((P2_P1_P2_HOLD == 1'b0) & (P2_P1_P2_RequestPending == 1'b1))) begin
                            $display(";A 5085");		//(= (bv-and (bv-comp P2_P1_P2_HOLD  0b0) (bv-comp P2_P1_P2_RequestPending  0b1))   0b1)) ;5085
                            P2_P1_P2_State <= #1 3'sb010; $display(";A 5087");		//(= P2_P1_P2_State    0b010)) ;5087
                        end
                        else begin
                            $display(";A 5086");		//(= (bv-and (bv-comp P2_P1_P2_HOLD  0b0) (bv-comp P2_P1_P2_RequestPending  0b1))   0b0)) ;5086
                            if (((P2_P1_P2_HOLD == 1'b0) & (P2_P1_P2_RequestPending == 1'b0))) begin
                                $display(";A 5088");		//(= (bv-and (bv-comp P2_P1_P2_HOLD  0b0) (bv-comp P2_P1_P2_RequestPending  0b0))   0b1)) ;5088
                                P2_P1_P2_State <= #1 3'sb001; $display(";A 5090");		//(= P2_P1_P2_State    0b001)) ;5090
                            end
                            else begin
                                $display(";A 5089");		//(= (bv-and (bv-comp P2_P1_P2_HOLD  0b0) (bv-comp P2_P1_P2_RequestPending  0b0))   0b0)) ;5089
                                P2_P1_P2_State <= #1 3'sb101; $display(";A 5091");		//(= P2_P1_P2_State    0b101)) ;5091
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 5092");		//(= P2_P1_P2_State    0b110)) ;5092
                        P2_P1_P2_Address <= #1 ((P2_P1_P2_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 5093");		//(= P2_P1_P2_Address    (bv-smod (bv-sdiv P2_P1_P2_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;5093
                        P2_P1_P2_BE_n <= #1 P2_P1_P2_ByteEnable; $display(";A 5094");		//(= P2_P1_P2_BE_n    P2_P1_P2_ByteEnable )) ;5094
                        P2_P1_P2_M_IO_n <= #1 P2_P1_P2_MemoryFetch; $display(";A 5095");		//(= P2_P1_P2_M_IO_n    P2_P1_P2_MemoryFetch )) ;5095
                        if ((P2_P1_P2_ReadRequest == 1'b1)) begin
                            $display(";A 5096");		//(= (bv-comp P2_P1_P2_ReadRequest  0b1)   0b1)) ;5096
                            P2_P1_P2_W_R_n <= #1 1'b0; $display(";A 5098");		//(= P2_P1_P2_W_R_n    0b0)) ;5098
                        end
                        else begin
                            $display(";A 5097");		//(= (bv-comp P2_P1_P2_ReadRequest  0b1)   0b0)) ;5097
                            P2_P1_P2_W_R_n <= #1 1'b1; $display(";A 5099");		//(= P2_P1_P2_W_R_n    0b1)) ;5099
                        end
                        if ((P2_P1_P2_CodeFetch == 1'b1)) begin
                            $display(";A 5100");		//(= (bv-comp P2_P1_P2_CodeFetch  0b1)   0b1)) ;5100
                            P2_P1_P2_D_C_n <= #1 1'b0; $display(";A 5102");		//(= P2_P1_P2_D_C_n    0b0)) ;5102
                        end
                        else begin
                            $display(";A 5101");		//(= (bv-comp P2_P1_P2_CodeFetch  0b1)   0b0)) ;5101
                            P2_P1_P2_D_C_n <= #1 1'b1; $display(";A 5103");		//(= P2_P1_P2_D_C_n    0b1)) ;5103
                        end
                        P2_P1_P2_ADS_n <= #1 1'b0; $display(";A 5104");		//(= P2_P1_P2_ADS_n    0b0)) ;5104
                        if ((P2_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 5105");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5105
                            P2_P1_P2_State <= #1 3'sb100; $display(";A 5107");		//(= P2_P1_P2_State    0b100)) ;5107
                        end
                        else begin
                            $display(";A 5106");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5106
                            P2_P1_P2_State <= #1 3'sb110; $display(";A 5108");		//(= P2_P1_P2_State    0b110)) ;5108
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 5109");		//(= P2_P1_P2_State    0b111)) ;5109
                        if ((((P2_P1_P2_READY_n == 1'b1) & (P2_P1_P2_RequestPending == 1'b1)) & (P2_P1_P2_HOLD == 1'b0))) begin
                            $display(";A 5110");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b1) (bv-comp P2_P1_P2_RequestPending  0b1)) (bv-comp P2_P1_P2_HOLD  0b0))   0b1)) ;5110
                            P2_P1_P2_State <= #1 3'sb110; $display(";A 5112");		//(= P2_P1_P2_State    0b110)) ;5112
                        end
                        else begin
                            $display(";A 5111");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b1) (bv-comp P2_P1_P2_RequestPending  0b1)) (bv-comp P2_P1_P2_HOLD  0b0))   0b0)) ;5111
                            if (((P2_P1_P2_READY_n == 1'b0) & (P2_P1_P2_HOLD == 1'b1))) begin
                                $display(";A 5113");		//(= (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b1))   0b1)) ;5113
                                P2_P1_P2_State <= #1 3'sb101; $display(";A 5115");		//(= P2_P1_P2_State    0b101)) ;5115
                            end
                            else begin
                                $display(";A 5114");		//(= (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b1))   0b0)) ;5114
                                if ((((P2_P1_P2_READY_n == 1'b0) & (P2_P1_P2_HOLD == 1'b0)) & (P2_P1_P2_RequestPending == 1'b1))) begin
                                    $display(";A 5116");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b1))   0b1)) ;5116
                                    P2_P1_P2_State <= #1 3'sb010; $display(";A 5118");		//(= P2_P1_P2_State    0b010)) ;5118
                                end
                                else begin
                                    $display(";A 5117");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b1))   0b0)) ;5117
                                    if ((((P2_P1_P2_READY_n == 1'b0) & (P2_P1_P2_HOLD == 1'b0)) & (P2_P1_P2_RequestPending == 1'b0))) begin
                                        $display(";A 5119");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b0))   0b1)) ;5119
                                        P2_P1_P2_State <= #1 3'sb001; $display(";A 5121");		//(= P2_P1_P2_State    0b001)) ;5121
                                    end
                                    else begin
                                        $display(";A 5120");		//(= (bv-and (bv-and (bv-comp P2_P1_P2_READY_n  0b0) (bv-comp P2_P1_P2_HOLD  0b0)) (bv-comp P2_P1_P2_RequestPending  0b0))   0b0)) ;5120
                                        P2_P1_P2_State <= #1 3'sb111; $display(";A 5122");		//(= P2_P1_P2_State    0b111)) ;5122
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:7806
    always @(posedge P2_P1_P2_RESET or posedge P2_P1_P2_CLOCK) begin
        if ((P2_P1_P2_RESET == 1'b1)) begin
            $display(";A 5123");		//(= (bv-comp P2_P1_P2_RESET  0b1)   0b1)) ;5123
            P2_P1_P2_State2 = 4'sb0000; $display(";A 5125");		//(= P2_P1_P2_State2    0b0000)) ;5125
            P2_P1_P2_InstQueue[0] = 8'b00000000; $display(";A 5126");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5126
            P2_P1_P2_InstQueue[1] = 8'b00000000; $display(";A 5127");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5127
            P2_P1_P2_InstQueue[2] = 8'b00000000; $display(";A 5128");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5128
            P2_P1_P2_InstQueue[3] = 8'b00000000; $display(";A 5129");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5129
            P2_P1_P2_InstQueue[4] = 8'b00000000; $display(";A 5130");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5130
            P2_P1_P2_InstQueue[5] = 8'b00000000; $display(";A 5131");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5131
            P2_P1_P2_InstQueue[6] = 8'b00000000; $display(";A 5132");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5132
            P2_P1_P2_InstQueue[7] = 8'b00000000; $display(";A 5133");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5133
            P2_P1_P2_InstQueue[8] = 8'b00000000; $display(";A 5134");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5134
            P2_P1_P2_InstQueue[9] = 8'b00000000; $display(";A 5135");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5135
            P2_P1_P2_InstQueue[10] = 8'b00000000; $display(";A 5136");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5136
            P2_P1_P2_InstQueue[11] = 8'b00000000; $display(";A 5137");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5137
            P2_P1_P2_InstQueue[12] = 8'b00000000; $display(";A 5138");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5138
            P2_P1_P2_InstQueue[13] = 8'b00000000; $display(";A 5139");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5139
            P2_P1_P2_InstQueue[14] = 8'b00000000; $display(";A 5140");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5140
            P2_P1_P2_InstQueue[15] = 8'b00000000; $display(";A 5141");		//(= P2_P1_P2_InstQueue    0b00000000)) ;5141
            P2_P1_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 5142");		//(= P2_P1_P2_InstQueueRd_Addr    0b00000)) ;5142
            P2_P1_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 5143");		//(= P2_P1_P2_InstQueueWr_Addr    0b00000)) ;5143
            P2_P1_P2_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 5144");		//(= P2_P1_P2_InstAddrPointer    0b00000000000000000000000000000000)) ;5144
            P2_P1_P2_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 5145");		//(= P2_P1_P2_PhyAddrPointer    0b00000000000000000000000000000000)) ;5145
            P2_P1_P2_Extended = 1'b0; $display(";A 5146");		//(= P2_P1_P2_Extended    0b0)) ;5146
            P2_P1_P2_More = 1'b0; $display(";A 5147");		//(= P2_P1_P2_More    0b0)) ;5147
            P2_P1_P2_Flush = 1'b0; $display(";A 5148");		//(= P2_P1_P2_Flush    0b0)) ;5148
            P2_P1_P2_lWord = 16'sb0000000000000000; $display(";A 5149");		//(= P2_P1_P2_lWord    0b0000000000000000)) ;5149
            P2_P1_P2_uWord = 15'sb000000000000000; $display(";A 5150");		//(= P2_P1_P2_uWord    0b000000000000000)) ;5150
            P2_P1_P2_fWord = 32'sb00000000000000000000000000000000; $display(";A 5151");		//(= P2_P1_P2_fWord    0b00000000000000000000000000000000)) ;5151
            P2_P1_P2_CodeFetch <= #1 1'b0; $display(";A 5152");		//(= P2_P1_P2_CodeFetch    0b0)) ;5152
            P2_P1_P2_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 5153");		//(= P2_P1_P2_Datao    0b00000000000000000000000000000000)) ;5153
            P2_P1_P2_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 5154");		//(= P2_P1_P2_EAX    0b00000000000000000000000000000000)) ;5154
            P2_P1_P2_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 5155");		//(= P2_P1_P2_EBX    0b00000000000000000000000000000000)) ;5155
            P2_P1_P2_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 5156");		//(= P2_P1_P2_rEIP    0b00000000000000000000000000000000)) ;5156
            P2_P1_P2_ReadRequest <= #1 1'b0; $display(";A 5157");		//(= P2_P1_P2_ReadRequest    0b0)) ;5157
            P2_P1_P2_MemoryFetch <= #1 1'b0; $display(";A 5158");		//(= P2_P1_P2_MemoryFetch    0b0)) ;5158
            P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5159");		//(= P2_P1_P2_RequestPending    0b0)) ;5159
        end
        else begin
            $display(";A 5124");		//(= (bv-comp P2_P1_P2_RESET  0b1)   0b0)) ;5124
            case (P2_P1_P2_State2)
                4'b0000 :
                    begin
                        $display(";A 5160");		//(= P2_P1_P2_State2    0b0000)) ;5160
                        P2_P1_P2_PhyAddrPointer = P2_P1_P2_rEIP; $display(";A 5161");		//(= P2_P1_P2_PhyAddrPointer    P2_P1_P2_rEIP )) ;5161
                        P2_P1_P2_InstAddrPointer = P2_P1_P2_PhyAddrPointer; $display(";A 5162");		//(= P2_P1_P2_InstAddrPointer    P2_P1_P2_PhyAddrPointer )) ;5162
                        P2_P1_P2_State2 = 4'sb0001; $display(";A 5163");		//(= P2_P1_P2_State2    0b0001)) ;5163
                        P2_P1_P2_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 5164");		//(= P2_P1_P2_rEIP    0b00000000000011111111111111110000)) ;5164
                        P2_P1_P2_ReadRequest <= #1 1'b1; $display(";A 5165");		//(= P2_P1_P2_ReadRequest    0b1)) ;5165
                        P2_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 5166");		//(= P2_P1_P2_MemoryFetch    0b1)) ;5166
                        P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5167");		//(= P2_P1_P2_RequestPending    0b1)) ;5167
                    end
                4'b0001 :
                    begin
                        $display(";A 5168");		//(= P2_P1_P2_State2    0b0001)) ;5168
                        P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5169");		//(= P2_P1_P2_RequestPending    0b1)) ;5169
                        P2_P1_P2_ReadRequest <= #1 1'b1; $display(";A 5170");		//(= P2_P1_P2_ReadRequest    0b1)) ;5170
                        P2_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 5171");		//(= P2_P1_P2_MemoryFetch    0b1)) ;5171
                        P2_P1_P2_CodeFetch <= #1 1'b1; $display(";A 5172");		//(= P2_P1_P2_CodeFetch    0b1)) ;5172
                        if ((P2_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 5173");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5173
                            P2_P1_P2_State2 = 4'sb0010; $display(";A 5175");		//(= P2_P1_P2_State2    0b0010)) ;5175
                        end
                        else begin
                            $display(";A 5174");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5174
                            P2_P1_P2_State2 = 4'sb0001; $display(";A 5176");		//(= P2_P1_P2_State2    0b0001)) ;5176
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 5177");		//(= P2_P1_P2_State2    0b0010)) ;5177
                        P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5178");		//(= P2_P1_P2_RequestPending    0b0)) ;5178
                        P2_P1_P2_InstQueue[P2_P1_P2_InstQueueWr_Addr] = (P2_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 5179");		//(= P2_P1_P2_InstQueue    (bv-smod P2_P1_P2_Datai  0b00000000000000000000000100000000))) ;5179
                        P2_P1_P2_InstQueueWr_Addr = ((P2_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5180");		//(= P2_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5180
                        P2_P1_P2_InstQueue[P2_P1_P2_InstQueueWr_Addr] = (P2_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 5181");		//(= P2_P1_P2_InstQueue    (bv-smod P2_P1_P2_Datai  0b00000000000000000000000100000000))) ;5181
                        P2_P1_P2_InstQueueWr_Addr = ((P2_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5182");		//(= P2_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5182
                        if ((P2_P1_P2_StateBS16 == 1'b1)) begin
                            $display(";A 5183");		//(= (bv-comp P2_P1_P2_StateBS16  0b1)   0b1)) ;5183
                            P2_P1_P2_InstQueue[P2_P1_P2_InstQueueWr_Addr] = ((P2_P1_P2_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 5185");		//(= P2_P1_P2_InstQueue    (bv-smod (bv-sdiv P2_P1_P2_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;5185
                            P2_P1_P2_InstQueueWr_Addr = ((P2_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5186");		//(= P2_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5186
                            P2_P1_P2_InstQueue[P2_P1_P2_InstQueueWr_Addr] = ((P2_P1_P2_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 5187");		//(= P2_P1_P2_InstQueue    (bv-smod (bv-sdiv P2_P1_P2_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;5187
                            P2_P1_P2_InstQueueWr_Addr = ((P2_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5188");		//(= P2_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5188
                            P2_P1_P2_PhyAddrPointer = (P2_P1_P2_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 5189");		//(= P2_P1_P2_PhyAddrPointer    (bv-add P2_P1_P2_PhyAddrPointer  0b00000000000000000000000000000100))) ;5189
                            P2_P1_P2_State2 = 4'sb0101; $display(";A 5190");		//(= P2_P1_P2_State2    0b0101)) ;5190
                        end
                        else begin
                            $display(";A 5184");		//(= (bv-comp P2_P1_P2_StateBS16  0b1)   0b0)) ;5184
                            P2_P1_P2_PhyAddrPointer = (P2_P1_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5191");		//(= P2_P1_P2_PhyAddrPointer    (bv-add P2_P1_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;5191
                            if ((P2_P1_P2_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 5192");		//(= (bool-to-bv (bv-slt P2_P1_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;5192
                                P2_P1_P2_rEIP <= #1 (-P2_P1_P2_PhyAddrPointer); $display(";A 5194");		//(= P2_P1_P2_rEIP    (bv-neg P2_P1_P2_PhyAddrPointer ))) ;5194
                            end
                            else begin
                                $display(";A 5193");		//(= (bool-to-bv (bv-slt P2_P1_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;5193
                                P2_P1_P2_rEIP <= #1 P2_P1_P2_PhyAddrPointer; $display(";A 5195");		//(= P2_P1_P2_rEIP    P2_P1_P2_PhyAddrPointer )) ;5195
                            end
                            P2_P1_P2_State2 = 4'sb0011; $display(";A 5196");		//(= P2_P1_P2_State2    0b0011)) ;5196
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 5197");		//(= P2_P1_P2_State2    0b0011)) ;5197
                        P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5198");		//(= P2_P1_P2_RequestPending    0b1)) ;5198
                        if ((P2_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 5199");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5199
                            P2_P1_P2_State2 = 4'sb0100; $display(";A 5201");		//(= P2_P1_P2_State2    0b0100)) ;5201
                        end
                        else begin
                            $display(";A 5200");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5200
                            P2_P1_P2_State2 = 4'sb0011; $display(";A 5202");		//(= P2_P1_P2_State2    0b0011)) ;5202
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 5203");		//(= P2_P1_P2_State2    0b0100)) ;5203
                        P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5204");		//(= P2_P1_P2_RequestPending    0b0)) ;5204
                        P2_P1_P2_InstQueue[P2_P1_P2_InstQueueWr_Addr] = (P2_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 5205");		//(= P2_P1_P2_InstQueue    (bv-smod P2_P1_P2_Datai  0b00000000000000000000000100000000))) ;5205
                        P2_P1_P2_InstQueueWr_Addr = ((P2_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5206");		//(= P2_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5206
                        P2_P1_P2_InstQueue[P2_P1_P2_InstQueueWr_Addr] = (P2_P1_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 5207");		//(= P2_P1_P2_InstQueue    (bv-smod P2_P1_P2_Datai  0b00000000000000000000000100000000))) ;5207
                        P2_P1_P2_InstQueueWr_Addr = ((P2_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5208");		//(= P2_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5208
                        P2_P1_P2_PhyAddrPointer = (P2_P1_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5209");		//(= P2_P1_P2_PhyAddrPointer    (bv-add P2_P1_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;5209
                        P2_P1_P2_State2 = 4'sb0101; $display(";A 5210");		//(= P2_P1_P2_State2    0b0101)) ;5210
                    end
                4'b0101 :
                    begin
                        $display(";A 5211");		//(= P2_P1_P2_State2    0b0101)) ;5211
                        case (P2_P1_P2_InstQueue[P2_P1_P2_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 5212");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b10010000)) ;5212
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5213");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5213
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5214");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5214
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5215");		//(= P2_P1_P2_Flush    0b0)) ;5215
                                    P2_P1_P2_More = 1'b0; $display(";A 5216");		//(= P2_P1_P2_More    0b0)) ;5216
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 5217");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b01100110)) ;5217
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5218");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5218
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5219");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5219
                                    P2_P1_P2_Extended = 1'b1; $display(";A 5220");		//(= P2_P1_P2_Extended    0b1)) ;5220
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5221");		//(= P2_P1_P2_Flush    0b0)) ;5221
                                    P2_P1_P2_More = 1'b0; $display(";A 5222");		//(= P2_P1_P2_More    0b0)) ;5222
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 5223");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b11101011)) ;5223
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 5224");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;5224
                                        if ((P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 5226");		//(= (bool-to-bv (bv-gt P2_P1_P2_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;5226
                                            P2_P1_P2_PhyAddrPointer = ((P2_P1_P2_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 5228");		//(= P2_P1_P2_PhyAddrPointer    (bv-sub (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P2_P1_P2_InstQueue 0 )))) ;5228
                                            P2_P1_P2_InstAddrPointer = P2_P1_P2_PhyAddrPointer; $display(";A 5229");		//(= P2_P1_P2_InstAddrPointer    P2_P1_P2_PhyAddrPointer )) ;5229
                                        end
                                        else begin
                                            $display(";A 5227");		//(= (bool-to-bv (bv-gt P2_P1_P2_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;5227
                                            P2_P1_P2_PhyAddrPointer = ((P2_P1_P2_InstAddrPointer + 32'b00000000000000000000000000000010) + P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 5230");		//(= P2_P1_P2_PhyAddrPointer    (bv-add (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000010) P2_P1_P2_InstQueue 0 ))) ;5230
                                            P2_P1_P2_InstAddrPointer = P2_P1_P2_PhyAddrPointer; $display(";A 5231");		//(= P2_P1_P2_InstAddrPointer    P2_P1_P2_PhyAddrPointer )) ;5231
                                        end
                                        P2_P1_P2_Flush = 1'b1; $display(";A 5232");		//(= P2_P1_P2_Flush    0b1)) ;5232
                                        P2_P1_P2_More = 1'b0; $display(";A 5233");		//(= P2_P1_P2_More    0b0)) ;5233
                                    end
                                    else begin
                                        $display(";A 5225");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;5225
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5234");		//(= P2_P1_P2_Flush    0b0)) ;5234
                                        P2_P1_P2_More = 1'b1; $display(";A 5235");		//(= P2_P1_P2_More    0b1)) ;5235
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 5236");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b11101001)) ;5236
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 5237");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;5237
                                        P2_P1_P2_PhyAddrPointer = ((P2_P1_P2_InstAddrPointer + 32'b00000000000000000000000000000101) + P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 5239");		//(= P2_P1_P2_PhyAddrPointer    (bv-add (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000101) P2_P1_P2_InstQueue 0 ))) ;5239
                                        P2_P1_P2_InstAddrPointer = P2_P1_P2_PhyAddrPointer; $display(";A 5240");		//(= P2_P1_P2_InstAddrPointer    P2_P1_P2_PhyAddrPointer )) ;5240
                                        P2_P1_P2_Flush = 1'b1; $display(";A 5241");		//(= P2_P1_P2_Flush    0b1)) ;5241
                                        P2_P1_P2_More = 1'b0; $display(";A 5242");		//(= P2_P1_P2_More    0b0)) ;5242
                                    end
                                    else begin
                                        $display(";A 5238");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;5238
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5243");		//(= P2_P1_P2_Flush    0b0)) ;5243
                                        P2_P1_P2_More = 1'b1; $display(";A 5244");		//(= P2_P1_P2_More    0b1)) ;5244
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 5245");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b11101010)) ;5245
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5246");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5246
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5247");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5247
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5248");		//(= P2_P1_P2_Flush    0b0)) ;5248
                                    P2_P1_P2_More = 1'b0; $display(";A 5249");		//(= P2_P1_P2_More    0b0)) ;5249
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 5250");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b10110000)) ;5250
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5251");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5251
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5252");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5252
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5253");		//(= P2_P1_P2_Flush    0b0)) ;5253
                                    P2_P1_P2_More = 1'b0; $display(";A 5254");		//(= P2_P1_P2_More    0b0)) ;5254
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 5255");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b10111000)) ;5255
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 5256");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;5256
                                        P2_P1_P2_EAX <= #1 ((((P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 5258");		//(= P2_P1_P2_EAX    (bv-add (bv-add (bv-add (bv-mul P2_P1_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P1_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P1_P2_InstQueue 0  0b00000000000000000000000100000000)) P2_P1_P2_InstQueue 0 ))) ;5258
                                        P2_P1_P2_More = 1'b0; $display(";A 5259");		//(= P2_P1_P2_More    0b0)) ;5259
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5260");		//(= P2_P1_P2_Flush    0b0)) ;5260
                                        P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 5261");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;5261
                                        P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 5262");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;5262
                                    end
                                    else begin
                                        $display(";A 5257");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;5257
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5263");		//(= P2_P1_P2_Flush    0b0)) ;5263
                                        P2_P1_P2_More = 1'b1; $display(";A 5264");		//(= P2_P1_P2_More    0b1)) ;5264
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 5265");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b10111011)) ;5265
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 5266");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;5266
                                        P2_P1_P2_EBX <= #1 ((((P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P1_P2_InstQueue[((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 5268");		//(= P2_P1_P2_EBX    (bv-add (bv-add (bv-add (bv-mul P2_P1_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P1_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P1_P2_InstQueue 0  0b00000000000000000000000100000000)) P2_P1_P2_InstQueue 0 ))) ;5268
                                        P2_P1_P2_More = 1'b0; $display(";A 5269");		//(= P2_P1_P2_More    0b0)) ;5269
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5270");		//(= P2_P1_P2_Flush    0b0)) ;5270
                                        P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 5271");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;5271
                                        P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 5272");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;5272
                                    end
                                    else begin
                                        $display(";A 5267");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;5267
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5273");		//(= P2_P1_P2_Flush    0b0)) ;5273
                                        P2_P1_P2_More = 1'b1; $display(";A 5274");		//(= P2_P1_P2_More    0b1)) ;5274
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 5275");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b10001011)) ;5275
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5276");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5276
                                        if ((P2_P1_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 5278");		//(= (bool-to-bv (bv-slt P2_P1_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;5278
                                            P2_P1_P2_rEIP <= #1 (-P2_P1_P2_EBX); $display(";A 5280");		//(= P2_P1_P2_rEIP    (bv-neg P2_P1_P2_EBX ))) ;5280
                                        end
                                        else begin
                                            $display(";A 5279");		//(= (bool-to-bv (bv-slt P2_P1_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;5279
                                            P2_P1_P2_rEIP <= #1 P2_P1_P2_EBX; $display(";A 5281");		//(= P2_P1_P2_rEIP    P2_P1_P2_EBX )) ;5281
                                        end
                                        P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5282");		//(= P2_P1_P2_RequestPending    0b1)) ;5282
                                        P2_P1_P2_ReadRequest <= #1 1'b1; $display(";A 5283");		//(= P2_P1_P2_ReadRequest    0b1)) ;5283
                                        P2_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 5284");		//(= P2_P1_P2_MemoryFetch    0b1)) ;5284
                                        P2_P1_P2_CodeFetch <= #1 1'b0; $display(";A 5285");		//(= P2_P1_P2_CodeFetch    0b0)) ;5285
                                        if ((P2_P1_P2_READY_n == 1'b0)) begin
                                            $display(";A 5286");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5286
                                            P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5288");		//(= P2_P1_P2_RequestPending    0b0)) ;5288
                                            P2_P1_P2_uWord = (P2_P1_P2_Datai % 32'b00000000000000001000000000000000); $display(";A 5289");		//(= P2_P1_P2_uWord    (bv-smod P2_P1_P2_Datai  0b00000000000000001000000000000000))) ;5289
                                            if ((P2_P1_P2_StateBS16 == 1'b1)) begin
                                                $display(";A 5290");		//(= (bv-comp P2_P1_P2_StateBS16  0b1)   0b1)) ;5290
                                                P2_P1_P2_lWord = (P2_P1_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 5292");		//(= P2_P1_P2_lWord    (bv-smod P2_P1_P2_Datai  0b00000000000000010000000000000000))) ;5292
                                            end
                                            else begin
                                                $display(";A 5291");		//(= (bv-comp P2_P1_P2_StateBS16  0b1)   0b0)) ;5291
                                                P2_P1_P2_rEIP <= #1 (P2_P1_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 5293");		//(= P2_P1_P2_rEIP    (bv-add P2_P1_P2_rEIP  0b00000000000000000000000000000010))) ;5293
                                                P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5294");		//(= P2_P1_P2_RequestPending    0b1)) ;5294
                                                if ((P2_P1_P2_READY_n == 1'b0)) begin
                                                    $display(";A 5295");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5295
                                                    P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5297");		//(= P2_P1_P2_RequestPending    0b0)) ;5297
                                                    P2_P1_P2_lWord = (P2_P1_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 5298");		//(= P2_P1_P2_lWord    (bv-smod P2_P1_P2_Datai  0b00000000000000010000000000000000))) ;5298
                                                end
                                                else begin
                                                    $display(";A 5296");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5296
                                                end
                                            end
                                            if ((P2_P1_P2_READY_n == 1'b0)) begin
                                                $display(";A 5299");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5299
                                                P2_P1_P2_EAX <= #1 ((P2_P1_P2_uWord * 32'b00000000000000010000000000000000) + P2_P1_P2_lWord); $display(";A 5301");		//(= P2_P1_P2_EAX    (bv-add (bv-mul P2_P1_P2_uWord  0b00000000000000010000000000000000) P2_P1_P2_lWord ))) ;5301
                                                P2_P1_P2_More = 1'b0; $display(";A 5302");		//(= P2_P1_P2_More    0b0)) ;5302
                                                P2_P1_P2_Flush = 1'b0; $display(";A 5303");		//(= P2_P1_P2_Flush    0b0)) ;5303
                                                P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5304");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;5304
                                                P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5305");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5305
                                            end
                                            else begin
                                                $display(";A 5300");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5300
                                            end
                                        end
                                        else begin
                                            $display(";A 5287");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5287
                                        end
                                    end
                                    else begin
                                        $display(";A 5277");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5277
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5306");		//(= P2_P1_P2_Flush    0b0)) ;5306
                                        P2_P1_P2_More = 1'b1; $display(";A 5307");		//(= P2_P1_P2_More    0b1)) ;5307
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 5308");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b10001001)) ;5308
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5309");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5309
                                        if ((P2_P1_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 5311");		//(= (bool-to-bv (bv-slt P2_P1_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;5311
                                            P2_P1_P2_rEIP <= #1 P2_P1_P2_EBX; $display(";A 5313");		//(= P2_P1_P2_rEIP    P2_P1_P2_EBX )) ;5313
                                        end
                                        else begin
                                            $display(";A 5312");		//(= (bool-to-bv (bv-slt P2_P1_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;5312
                                            P2_P1_P2_rEIP <= #1 P2_P1_P2_EBX; $display(";A 5314");		//(= P2_P1_P2_rEIP    P2_P1_P2_EBX )) ;5314
                                        end
                                        P2_P1_P2_lWord = (P2_P1_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 5315");		//(= P2_P1_P2_lWord    (bv-smod P2_P1_P2_EAX  0b00000000000000010000000000000000))) ;5315
                                        P2_P1_P2_uWord = ((P2_P1_P2_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 5316");		//(= P2_P1_P2_uWord    (bv-smod (bv-sdiv P2_P1_P2_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;5316
                                        P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5317");		//(= P2_P1_P2_RequestPending    0b1)) ;5317
                                        P2_P1_P2_ReadRequest <= #1 1'b0; $display(";A 5318");		//(= P2_P1_P2_ReadRequest    0b0)) ;5318
                                        P2_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 5319");		//(= P2_P1_P2_MemoryFetch    0b1)) ;5319
                                        P2_P1_P2_CodeFetch <= #1 1'b0; $display(";A 5320");		//(= P2_P1_P2_CodeFetch    0b0)) ;5320
                                        if (((P2_P1_P2_State == 32'b00000000000000000000000000000010) | (P2_P1_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 5321");		//(= (bv-or (bv-comp P2_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P2_State  0b00000000000000000000000000000100))   0b1)) ;5321
                                            P2_P1_P2_Datao <= #1 ((P2_P1_P2_uWord * 32'b00000000000000010000000000000000) + P2_P1_P2_lWord); $display(";A 5323");		//(= P2_P1_P2_Datao    (bv-add (bv-mul P2_P1_P2_uWord  0b00000000000000010000000000000000) P2_P1_P2_lWord ))) ;5323
                                            if ((P2_P1_P2_READY_n == 1'b0)) begin
                                                $display(";A 5324");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5324
                                                P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5326");		//(= P2_P1_P2_RequestPending    0b0)) ;5326
                                                if ((P2_P1_P2_StateBS16 == 1'b0)) begin
                                                    $display(";A 5327");		//(= (bv-comp P2_P1_P2_StateBS16  0b0)   0b1)) ;5327
                                                    P2_P1_P2_rEIP <= #1 (P2_P1_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 5329");		//(= P2_P1_P2_rEIP    (bv-add P2_P1_P2_rEIP  0b00000000000000000000000000000010))) ;5329
                                                    P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5330");		//(= P2_P1_P2_RequestPending    0b1)) ;5330
                                                    P2_P1_P2_ReadRequest <= #1 1'b0; $display(";A 5331");		//(= P2_P1_P2_ReadRequest    0b0)) ;5331
                                                    P2_P1_P2_MemoryFetch <= #1 1'b1; $display(";A 5332");		//(= P2_P1_P2_MemoryFetch    0b1)) ;5332
                                                    P2_P1_P2_CodeFetch <= #1 1'b0; $display(";A 5333");		//(= P2_P1_P2_CodeFetch    0b0)) ;5333
                                                    P2_P1_P2_State2 = 4'sb0110; $display(";A 5334");		//(= P2_P1_P2_State2    0b0110)) ;5334
                                                end
                                                else begin
                                                    $display(";A 5328");		//(= (bv-comp P2_P1_P2_StateBS16  0b0)   0b0)) ;5328
                                                end
                                                P2_P1_P2_More = 1'b0; $display(";A 5335");		//(= P2_P1_P2_More    0b0)) ;5335
                                                P2_P1_P2_Flush = 1'b0; $display(";A 5336");		//(= P2_P1_P2_Flush    0b0)) ;5336
                                                P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5337");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;5337
                                                P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5338");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5338
                                            end
                                            else begin
                                                $display(";A 5325");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5325
                                            end
                                        end
                                        else begin
                                            $display(";A 5322");		//(= (bv-or (bv-comp P2_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P2_State  0b00000000000000000000000000000100))   0b0)) ;5322
                                        end
                                    end
                                    else begin
                                        $display(";A 5310");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5310
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5339");		//(= P2_P1_P2_Flush    0b0)) ;5339
                                        P2_P1_P2_More = 1'b1; $display(";A 5340");		//(= P2_P1_P2_More    0b1)) ;5340
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 5341");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b11100100)) ;5341
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5342");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5342
                                        P2_P1_P2_rEIP <= #1 (P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 5344");		//(= P2_P1_P2_rEIP    (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;5344
                                        P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5345");		//(= P2_P1_P2_RequestPending    0b1)) ;5345
                                        P2_P1_P2_ReadRequest <= #1 1'b1; $display(";A 5346");		//(= P2_P1_P2_ReadRequest    0b1)) ;5346
                                        P2_P1_P2_MemoryFetch <= #1 1'b0; $display(";A 5347");		//(= P2_P1_P2_MemoryFetch    0b0)) ;5347
                                        P2_P1_P2_CodeFetch <= #1 1'b0; $display(";A 5348");		//(= P2_P1_P2_CodeFetch    0b0)) ;5348
                                        if ((P2_P1_P2_READY_n == 1'b0)) begin
                                            $display(";A 5349");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5349
                                            P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5351");		//(= P2_P1_P2_RequestPending    0b0)) ;5351
                                            P2_P1_P2_EAX <= #1 P2_P1_P2_Datai; $display(";A 5352");		//(= P2_P1_P2_EAX    P2_P1_P2_Datai )) ;5352
                                            P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5353");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;5353
                                            P2_P1_P2_InstQueueRd_Addr = (P2_P1_P2_InstQueueRd_Addr + 5'b00010); $display(";A 5354");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-add P2_P1_P2_InstQueueRd_Addr  0b00010))) ;5354
                                            P2_P1_P2_Flush = 1'b0; $display(";A 5355");		//(= P2_P1_P2_Flush    0b0)) ;5355
                                            P2_P1_P2_More = 1'b0; $display(";A 5356");		//(= P2_P1_P2_More    0b0)) ;5356
                                        end
                                        else begin
                                            $display(";A 5350");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5350
                                        end
                                    end
                                    else begin
                                        $display(";A 5343");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5343
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5357");		//(= P2_P1_P2_Flush    0b0)) ;5357
                                        P2_P1_P2_More = 1'b1; $display(";A 5358");		//(= P2_P1_P2_More    0b1)) ;5358
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 5359");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b11100110)) ;5359
                                    if (((P2_P1_P2_InstQueueWr_Addr - P2_P1_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5360");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5360
                                        P2_P1_P2_rEIP <= #1 (P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 5362");		//(= P2_P1_P2_rEIP    (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;5362
                                        P2_P1_P2_RequestPending <= #1 1'b1; $display(";A 5363");		//(= P2_P1_P2_RequestPending    0b1)) ;5363
                                        P2_P1_P2_ReadRequest <= #1 1'b0; $display(";A 5364");		//(= P2_P1_P2_ReadRequest    0b0)) ;5364
                                        P2_P1_P2_MemoryFetch <= #1 1'b0; $display(";A 5365");		//(= P2_P1_P2_MemoryFetch    0b0)) ;5365
                                        P2_P1_P2_CodeFetch <= #1 1'b0; $display(";A 5366");		//(= P2_P1_P2_CodeFetch    0b0)) ;5366
                                        if (((P2_P1_P2_State == 32'b00000000000000000000000000000010) | (P2_P1_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 5367");		//(= (bv-or (bv-comp P2_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P2_State  0b00000000000000000000000000000100))   0b1)) ;5367
                                            P2_P1_P2_fWord = (P2_P1_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 5369");		//(= P2_P1_P2_fWord    (bv-smod P2_P1_P2_EAX  0b00000000000000010000000000000000))) ;5369
                                            P2_P1_P2_Datao <= #1 P2_P1_P2_fWord; $display(";A 5370");		//(= P2_P1_P2_Datao    P2_P1_P2_fWord )) ;5370
                                            if ((P2_P1_P2_READY_n == 1'b0)) begin
                                                $display(";A 5371");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5371
                                                P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5373");		//(= P2_P1_P2_RequestPending    0b0)) ;5373
                                                P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5374");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;5374
                                                P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5375");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5375
                                                P2_P1_P2_Flush = 1'b0; $display(";A 5376");		//(= P2_P1_P2_Flush    0b0)) ;5376
                                                P2_P1_P2_More = 1'b0; $display(";A 5377");		//(= P2_P1_P2_More    0b0)) ;5377
                                            end
                                            else begin
                                                $display(";A 5372");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5372
                                            end
                                        end
                                        else begin
                                            $display(";A 5368");		//(= (bv-or (bv-comp P2_P1_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P2_State  0b00000000000000000000000000000100))   0b0)) ;5368
                                        end
                                    end
                                    else begin
                                        $display(";A 5361");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P2_InstQueueWr_Addr  P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5361
                                        P2_P1_P2_Flush = 1'b0; $display(";A 5378");		//(= P2_P1_P2_Flush    0b0)) ;5378
                                        P2_P1_P2_More = 1'b1; $display(";A 5379");		//(= P2_P1_P2_More    0b1)) ;5379
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 5380");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b00000100)) ;5380
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5381");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5381
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5382");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5382
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5383");		//(= P2_P1_P2_Flush    0b0)) ;5383
                                    P2_P1_P2_More = 1'b0; $display(";A 5384");		//(= P2_P1_P2_More    0b0)) ;5384
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 5385");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b00000101)) ;5385
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5386");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5386
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5387");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5387
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5388");		//(= P2_P1_P2_Flush    0b0)) ;5388
                                    P2_P1_P2_More = 1'b0; $display(";A 5389");		//(= P2_P1_P2_More    0b0)) ;5389
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 5390");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b11010000)) ;5390
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5391");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;5391
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5392");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5392
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5393");		//(= P2_P1_P2_Flush    0b0)) ;5393
                                    P2_P1_P2_More = 1'b0; $display(";A 5394");		//(= P2_P1_P2_More    0b0)) ;5394
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 5395");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b11000000)) ;5395
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5396");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;5396
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5397");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5397
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5398");		//(= P2_P1_P2_Flush    0b0)) ;5398
                                    P2_P1_P2_More = 1'b0; $display(";A 5399");		//(= P2_P1_P2_More    0b0)) ;5399
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 5400");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b01000000)) ;5400
                                    P2_P1_P2_EAX <= #1 (P2_P1_P2_EAX + 32'sb00000000000000000000000000000001); $display(";A 5401");		//(= P2_P1_P2_EAX    (bv-add P2_P1_P2_EAX  0b00000000000000000000000000000001))) ;5401
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5402");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5402
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5403");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5403
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5404");		//(= P2_P1_P2_Flush    0b0)) ;5404
                                    P2_P1_P2_More = 1'b0; $display(";A 5405");		//(= P2_P1_P2_More    0b0)) ;5405
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 5406");		//(= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr )   0b01000011)) ;5406
                                    P2_P1_P2_EBX <= #1 (P2_P1_P2_EBX + 32'sb00000000000000000000000000000001); $display(";A 5407");		//(= P2_P1_P2_EBX    (bv-add P2_P1_P2_EBX  0b00000000000000000000000000000001))) ;5407
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5408");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5408
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5409");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5409
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5410");		//(= P2_P1_P2_Flush    0b0)) ;5410
                                    P2_P1_P2_More = 1'b0; $display(";A 5411");		//(= P2_P1_P2_More    0b0)) ;5411
                                end
                            default:
                                begin
                                    $display(";A 5412");		//(= (and (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b10010000) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b01100110) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b11101011) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b11101001) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b11101010) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b10110000) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b10111000) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b10111011) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b10001011) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b10001001) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b11100100) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b11100110) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b00000100) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b00000101) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b11010000) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b11000000) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b01000000) (/= ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ) 0b01000011))   true)) ;5412
                                    P2_P1_P2_InstAddrPointer = (P2_P1_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5413");		//(= P2_P1_P2_InstAddrPointer    (bv-add P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;5413
                                    P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5414");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5414
                                    P2_P1_P2_Flush = 1'b0; $display(";A 5415");		//(= P2_P1_P2_Flush    0b0)) ;5415
                                    P2_P1_P2_More = 1'b0; $display(";A 5416");		//(= P2_P1_P2_More    0b0)) ;5416
                                end
                        endcase
                        if (((~(P2_P1_P2_InstQueueRd_Addr < P2_P1_P2_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P2_P1_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P2_P1_P2_Flush) | P2_P1_P2_More))) begin
                            $display(";A 5417");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P1_P2_InstQueueRd_Addr  P2_P1_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P1_P2_Flush ) P2_P1_P2_More ))   0b1)) ;5417
                            P2_P1_P2_State2 = 4'sb0111; $display(";A 5419");		//(= P2_P1_P2_State2    0b0111)) ;5419
                        end
                        else begin
                            $display(";A 5418");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P1_P2_InstQueueRd_Addr  P2_P1_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P1_P2_Flush ) P2_P1_P2_More ))   0b0)) ;5418
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 5420");		//(= P2_P1_P2_State2    0b0110)) ;5420
                        P2_P1_P2_Datao <= #1 ((P2_P1_P2_uWord * 32'b00000000000000010000000000000000) + P2_P1_P2_lWord); $display(";A 5421");		//(= P2_P1_P2_Datao    (bv-add (bv-mul P2_P1_P2_uWord  0b00000000000000010000000000000000) P2_P1_P2_lWord ))) ;5421
                        if ((P2_P1_P2_READY_n == 1'b0)) begin
                            $display(";A 5422");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b1)) ;5422
                            P2_P1_P2_RequestPending <= #1 1'b0; $display(";A 5424");		//(= P2_P1_P2_RequestPending    0b0)) ;5424
                            P2_P1_P2_State2 = 4'sb0101; $display(";A 5425");		//(= P2_P1_P2_State2    0b0101)) ;5425
                        end
                        else begin
                            $display(";A 5423");		//(= (bv-comp P2_P1_P2_READY_n  0b0)   0b0)) ;5423
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 5426");		//(= P2_P1_P2_State2    0b0111)) ;5426
                        if (P2_P1_P2_Flush) begin
                            $display(";A 5427");		//(= P2_P1_P2_Flush    0b1)) ;5427
                            P2_P1_P2_InstQueueRd_Addr = 5'sb00001; $display(";A 5429");		//(= P2_P1_P2_InstQueueRd_Addr    0b00001)) ;5429
                            P2_P1_P2_InstQueueWr_Addr = 5'sb00001; $display(";A 5430");		//(= P2_P1_P2_InstQueueWr_Addr    0b00001)) ;5430
                            if ((P2_P1_P2_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 5431");		//(= (bool-to-bv (bv-slt P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;5431
                                P2_P1_P2_fWord = (-P2_P1_P2_InstAddrPointer); $display(";A 5433");		//(= P2_P1_P2_fWord    (bv-neg P2_P1_P2_InstAddrPointer ))) ;5433
                            end
                            else begin
                                $display(";A 5432");		//(= (bool-to-bv (bv-slt P2_P1_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;5432
                                P2_P1_P2_fWord = P2_P1_P2_InstAddrPointer; $display(";A 5434");		//(= P2_P1_P2_fWord    P2_P1_P2_InstAddrPointer )) ;5434
                            end
                            if (((P2_P1_P2_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 5435");		//(= (bv-comp (bv-smod P2_P1_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;5435
                                P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + (P2_P1_P2_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 5437");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  (bv-smod P2_P1_P2_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;5437
                            end
                            else begin
                                $display(";A 5436");		//(= (bv-comp (bv-smod P2_P1_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;5436
                            end
                        end
                        else begin
                            $display(";A 5428");		//(= P2_P1_P2_Flush    0b0)) ;5428
                        end
                        if (((32'b00000000000000000000000000001111 - P2_P1_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 5438");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;5438
                            P2_P1_P2_State2 = 4'sb1000; $display(";A 5440");		//(= P2_P1_P2_State2    0b1000)) ;5440
                            P2_P1_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 5441");		//(= P2_P1_P2_InstQueueWr_Addr    0b00000)) ;5441
                        end
                        else begin
                            $display(";A 5439");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;5439
                            P2_P1_P2_State2 = 4'sb1001; $display(";A 5442");		//(= P2_P1_P2_State2    0b1001)) ;5442
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 5443");		//(= P2_P1_P2_State2    0b1000)) ;5443
                        if ((P2_P1_P2_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 5444");		//(= (bool-to-bv (bv-le P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;5444
                            P2_P1_P2_InstQueue[P2_P1_P2_InstQueueWr_Addr] = P2_P1_P2_InstQueue[P2_P1_P2_InstQueueRd_Addr]; $display(";A 5446");		//(= P2_P1_P2_InstQueue    ( P2_P1_P2_InstQueue P2_P1_P2_InstQueueRd_Addr ))) ;5446
                            P2_P1_P2_InstQueueRd_Addr = ((P2_P1_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5447");		//(= P2_P1_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5447
                            P2_P1_P2_InstQueueWr_Addr = ((P2_P1_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5448");		//(= P2_P1_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5448
                            P2_P1_P2_State2 = 4'sb1000; $display(";A 5449");		//(= P2_P1_P2_State2    0b1000)) ;5449
                        end
                        else begin
                            $display(";A 5445");		//(= (bool-to-bv (bv-le P2_P1_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;5445
                            P2_P1_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 5450");		//(= P2_P1_P2_InstQueueRd_Addr    0b00000)) ;5450
                            P2_P1_P2_State2 = 4'sb1001; $display(";A 5451");		//(= P2_P1_P2_State2    0b1001)) ;5451
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 5452");		//(= P2_P1_P2_State2    0b1001)) ;5452
                        P2_P1_P2_rEIP <= #1 P2_P1_P2_PhyAddrPointer; $display(";A 5453");		//(= P2_P1_P2_rEIP    P2_P1_P2_PhyAddrPointer )) ;5453
                        P2_P1_P2_State2 = 4'sb0001; $display(";A 5454");		//(= P2_P1_P2_State2    0b0001)) ;5454
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:8245
    always @(posedge P2_P1_P2_RESET or posedge P2_P1_P2_CLOCK) begin
        if ((P2_P1_P2_RESET == 1'b1)) begin
            $display(";A 5455");		//(= (bv-comp P2_P1_P2_RESET  0b1)   0b1)) ;5455
            P2_P1_P2_ByteEnable <= #1 4'b0000; $display(";A 5457");		//(= P2_P1_P2_ByteEnable    0b0000)) ;5457
            P2_P1_P2_NonAligned <= #1 1'b0; $display(";A 5458");		//(= P2_P1_P2_NonAligned    0b0)) ;5458
        end
        else begin
            $display(";A 5456");		//(= (bv-comp P2_P1_P2_RESET  0b1)   0b0)) ;5456
            case (P2_P1_P2_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 5459");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000000)) ;5459
                        case ((P2_P1_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 5460");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;5460
                                    P2_P1_P2_ByteEnable <= #1 4'b1110; $display(";A 5461");		//(= P2_P1_P2_ByteEnable    0b1110)) ;5461
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 5462");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;5462
                                    P2_P1_P2_ByteEnable <= #1 4'b1101; $display(";A 5463");		//(= P2_P1_P2_ByteEnable    0b1101)) ;5463
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 5464");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;5464
                                    P2_P1_P2_ByteEnable <= #1 4'b1011; $display(";A 5465");		//(= P2_P1_P2_ByteEnable    0b1011)) ;5465
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 5466");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;5466
                                    P2_P1_P2_ByteEnable <= #1 4'b0111; $display(";A 5467");		//(= P2_P1_P2_ByteEnable    0b0111)) ;5467
                                end
                            default:
                                begin
                                    $display(";A 5468");		//(= (and (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;5468
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 5469");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000001)) ;5469
                        case ((P2_P1_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 5470");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;5470
                                    P2_P1_P2_ByteEnable <= #1 4'b1100; $display(";A 5471");		//(= P2_P1_P2_ByteEnable    0b1100)) ;5471
                                    P2_P1_P2_NonAligned <= #1 1'b0; $display(";A 5472");		//(= P2_P1_P2_NonAligned    0b0)) ;5472
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 5473");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;5473
                                    P2_P1_P2_ByteEnable <= #1 4'b1001; $display(";A 5474");		//(= P2_P1_P2_ByteEnable    0b1001)) ;5474
                                    P2_P1_P2_NonAligned <= #1 1'b0; $display(";A 5475");		//(= P2_P1_P2_NonAligned    0b0)) ;5475
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 5476");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;5476
                                    P2_P1_P2_ByteEnable <= #1 4'b0011; $display(";A 5477");		//(= P2_P1_P2_ByteEnable    0b0011)) ;5477
                                    P2_P1_P2_NonAligned <= #1 1'b0; $display(";A 5478");		//(= P2_P1_P2_NonAligned    0b0)) ;5478
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 5479");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;5479
                                    P2_P1_P2_ByteEnable <= #1 4'b0111; $display(";A 5480");		//(= P2_P1_P2_ByteEnable    0b0111)) ;5480
                                    P2_P1_P2_NonAligned <= #1 1'b1; $display(";A 5481");		//(= P2_P1_P2_NonAligned    0b1)) ;5481
                                end
                            default:
                                begin
                                    $display(";A 5482");		//(= (and (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;5482
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 5483");		//(= P2_P1_P2_DataWidth    0b00000000000000000000000000000010)) ;5483
                        case ((P2_P1_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 5484");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;5484
                                    P2_P1_P2_ByteEnable <= #1 4'b0000; $display(";A 5485");		//(= P2_P1_P2_ByteEnable    0b0000)) ;5485
                                    P2_P1_P2_NonAligned <= #1 1'b0; $display(";A 5486");		//(= P2_P1_P2_NonAligned    0b0)) ;5486
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 5487");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;5487
                                    P2_P1_P2_ByteEnable <= #1 4'b0001; $display(";A 5488");		//(= P2_P1_P2_ByteEnable    0b0001)) ;5488
                                    P2_P1_P2_NonAligned <= #1 1'b1; $display(";A 5489");		//(= P2_P1_P2_NonAligned    0b1)) ;5489
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 5490");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;5490
                                    P2_P1_P2_NonAligned <= #1 1'b1; $display(";A 5491");		//(= P2_P1_P2_NonAligned    0b1)) ;5491
                                    P2_P1_P2_ByteEnable <= #1 4'b0011; $display(";A 5492");		//(= P2_P1_P2_ByteEnable    0b0011)) ;5492
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 5493");		//(= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;5493
                                    P2_P1_P2_NonAligned <= #1 1'b1; $display(";A 5494");		//(= P2_P1_P2_NonAligned    0b1)) ;5494
                                    P2_P1_P2_ByteEnable <= #1 4'b0111; $display(";A 5495");		//(= P2_P1_P2_ByteEnable    0b0111)) ;5495
                                end
                            default:
                                begin
                                    $display(";A 5496");		//(= (and (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;5496
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 5497");		//(= (and (/= P2_P1_P2_DataWidth  0b00000000000000000000000000000000) (/= P2_P1_P2_DataWidth  0b00000000000000000000000000000001) (/= P2_P1_P2_DataWidth  0b00000000000000000000000000000010))   true)) ;5497
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:8433
    always @(posedge P2_P1_P3_RESET or posedge P2_P1_P3_CLOCK) begin
        if ((P2_P1_P3_RESET == 1'b1)) begin
            $display(";A 5498");		//(= (bv-comp P2_P1_P3_RESET  0b1)   0b1)) ;5498
            P2_P1_P3_BE_n <= #1 4'b0000; $display(";A 5500");		//(= P2_P1_P3_BE_n    0b0000)) ;5500
            P2_P1_P3_Address <= #1 30'sb000000000000000000000000000000; $display(";A 5501");		//(= P2_P1_P3_Address    0b000000000000000000000000000000)) ;5501
            P2_P1_P3_W_R_n <= #1 1'b0; $display(";A 5502");		//(= P2_P1_P3_W_R_n    0b0)) ;5502
            P2_P1_P3_D_C_n <= #1 1'b0; $display(";A 5503");		//(= P2_P1_P3_D_C_n    0b0)) ;5503
            P2_P1_P3_M_IO_n <= #1 1'b0; $display(";A 5504");		//(= P2_P1_P3_M_IO_n    0b0)) ;5504
            P2_P1_P3_ADS_n <= #1 1'b0; $display(";A 5505");		//(= P2_P1_P3_ADS_n    0b0)) ;5505
            P2_P1_P3_State <= #1 3'sb000; $display(";A 5506");		//(= P2_P1_P3_State    0b000)) ;5506
            P2_P1_P3_StateNA <= #1 1'b0; $display(";A 5507");		//(= P2_P1_P3_StateNA    0b0)) ;5507
            P2_P1_P3_StateBS16 <= #1 1'b0; $display(";A 5508");		//(= P2_P1_P3_StateBS16    0b0)) ;5508
            P2_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 5509");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000000)) ;5509
        end
        else begin
            $display(";A 5499");		//(= (bv-comp P2_P1_P3_RESET  0b1)   0b0)) ;5499
            case (P2_P1_P3_State)
                3'b000 :
                    begin
                        $display(";A 5510");		//(= P2_P1_P3_State    0b000)) ;5510
                        P2_P1_P3_D_C_n <= #1 1'b1; $display(";A 5511");		//(= P2_P1_P3_D_C_n    0b1)) ;5511
                        P2_P1_P3_ADS_n <= #1 1'b1; $display(";A 5512");		//(= P2_P1_P3_ADS_n    0b1)) ;5512
                        P2_P1_P3_State <= #1 3'sb001; $display(";A 5513");		//(= P2_P1_P3_State    0b001)) ;5513
                        P2_P1_P3_StateNA <= #1 1'b1; $display(";A 5514");		//(= P2_P1_P3_StateNA    0b1)) ;5514
                        P2_P1_P3_StateBS16 <= #1 1'b1; $display(";A 5515");		//(= P2_P1_P3_StateBS16    0b1)) ;5515
                        P2_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 5516");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;5516
                        P2_P1_P3_State <= #1 3'sb001; $display(";A 5517");		//(= P2_P1_P3_State    0b001)) ;5517
                    end
                3'b001 :
                    begin
                        $display(";A 5518");		//(= P2_P1_P3_State    0b001)) ;5518
                        if ((P2_P1_P3_RequestPending == 1'b1)) begin
                            $display(";A 5519");		//(= (bv-comp P2_P1_P3_RequestPending  0b1)   0b1)) ;5519
                            P2_P1_P3_State <= #1 3'sb010; $display(";A 5521");		//(= P2_P1_P3_State    0b010)) ;5521
                        end
                        else begin
                            $display(";A 5520");		//(= (bv-comp P2_P1_P3_RequestPending  0b1)   0b0)) ;5520
                            if ((P2_P1_P3_HOLD == 1'b1)) begin
                                $display(";A 5522");		//(= (bv-comp P2_P1_P3_HOLD  0b1)   0b1)) ;5522
                                P2_P1_P3_State <= #1 3'sb101; $display(";A 5524");		//(= P2_P1_P3_State    0b101)) ;5524
                            end
                            else begin
                                $display(";A 5523");		//(= (bv-comp P2_P1_P3_HOLD  0b1)   0b0)) ;5523
                                P2_P1_P3_State <= #1 3'sb001; $display(";A 5525");		//(= P2_P1_P3_State    0b001)) ;5525
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 5526");		//(= P2_P1_P3_State    0b010)) ;5526
                        P2_P1_P3_Address <= #1 ((P2_P1_P3_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 5527");		//(= P2_P1_P3_Address    (bv-smod (bv-sdiv P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;5527
                        P2_P1_P3_BE_n <= #1 P2_P1_P3_ByteEnable; $display(";A 5528");		//(= P2_P1_P3_BE_n    P2_P1_P3_ByteEnable )) ;5528
                        P2_P1_P3_M_IO_n <= #1 P2_P1_P3_MemoryFetch; $display(";A 5529");		//(= P2_P1_P3_M_IO_n    P2_P1_P3_MemoryFetch )) ;5529
                        if ((P2_P1_P3_ReadRequest == 1'b1)) begin
                            $display(";A 5530");		//(= (bv-comp P2_P1_P3_ReadRequest  0b1)   0b1)) ;5530
                            P2_P1_P3_W_R_n <= #1 1'b0; $display(";A 5532");		//(= P2_P1_P3_W_R_n    0b0)) ;5532
                        end
                        else begin
                            $display(";A 5531");		//(= (bv-comp P2_P1_P3_ReadRequest  0b1)   0b0)) ;5531
                            P2_P1_P3_W_R_n <= #1 1'b1; $display(";A 5533");		//(= P2_P1_P3_W_R_n    0b1)) ;5533
                        end
                        if ((P2_P1_P3_CodeFetch == 1'b1)) begin
                            $display(";A 5534");		//(= (bv-comp P2_P1_P3_CodeFetch  0b1)   0b1)) ;5534
                            P2_P1_P3_D_C_n <= #1 1'b0; $display(";A 5536");		//(= P2_P1_P3_D_C_n    0b0)) ;5536
                        end
                        else begin
                            $display(";A 5535");		//(= (bv-comp P2_P1_P3_CodeFetch  0b1)   0b0)) ;5535
                            P2_P1_P3_D_C_n <= #1 1'b1; $display(";A 5537");		//(= P2_P1_P3_D_C_n    0b1)) ;5537
                        end
                        P2_P1_P3_ADS_n <= #1 1'b0; $display(";A 5538");		//(= P2_P1_P3_ADS_n    0b0)) ;5538
                        P2_P1_P3_State <= #1 3'sb011; $display(";A 5539");		//(= P2_P1_P3_State    0b011)) ;5539
                    end
                3'b011 :
                    begin
                        $display(";A 5540");		//(= P2_P1_P3_State    0b011)) ;5540
                        if ((((P2_P1_P3_READY_n == 1'b0) & (P2_P1_P3_HOLD == 1'b0)) & (P2_P1_P3_RequestPending == 1'b1))) begin
                            $display(";A 5541");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b1))   0b1)) ;5541
                            P2_P1_P3_State <= #1 3'sb010; $display(";A 5543");		//(= P2_P1_P3_State    0b010)) ;5543
                        end
                        else begin
                            $display(";A 5542");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b1))   0b0)) ;5542
                            if (((P2_P1_P3_READY_n == 1'b1) & (P2_P1_P3_NA_n == 1'b1))) begin
                                $display(";A 5544");		//(= (bv-and (bv-comp P2_P1_P3_READY_n  0b1) (bv-comp P2_P1_P3_NA_n  0b1))   0b1)) ;5544
                            end
                            else begin
                                $display(";A 5545");		//(= (bv-and (bv-comp P2_P1_P3_READY_n  0b1) (bv-comp P2_P1_P3_NA_n  0b1))   0b0)) ;5545
                                if ((((P2_P1_P3_RequestPending == 1'b1) | (P2_P1_P3_HOLD == 1'b1)) & ((P2_P1_P3_READY_n == 1'b1) & (P2_P1_P3_NA_n == 1'b0)))) begin
                                    $display(";A 5546");		//(= (bv-and (bv-or (bv-comp P2_P1_P3_RequestPending  0b1) (bv-comp P2_P1_P3_HOLD  0b1)) (bv-and (bv-comp P2_P1_P3_READY_n  0b1) (bv-comp P2_P1_P3_NA_n  0b0)))   0b1)) ;5546
                                    P2_P1_P3_State <= #1 3'sb111; $display(";A 5548");		//(= P2_P1_P3_State    0b111)) ;5548
                                end
                                else begin
                                    $display(";A 5547");		//(= (bv-and (bv-or (bv-comp P2_P1_P3_RequestPending  0b1) (bv-comp P2_P1_P3_HOLD  0b1)) (bv-and (bv-comp P2_P1_P3_READY_n  0b1) (bv-comp P2_P1_P3_NA_n  0b0)))   0b0)) ;5547
                                    if (((((P2_P1_P3_RequestPending == 1'b1) & (P2_P1_P3_HOLD == 1'b0)) & (P2_P1_P3_READY_n == 1'b1)) & (P2_P1_P3_NA_n == 1'b0))) begin
                                        $display(";A 5549");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P1_P3_RequestPending  0b1) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_READY_n  0b1)) (bv-comp P2_P1_P3_NA_n  0b0))   0b1)) ;5549
                                        P2_P1_P3_State <= #1 3'sb110; $display(";A 5551");		//(= P2_P1_P3_State    0b110)) ;5551
                                    end
                                    else begin
                                        $display(";A 5550");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P1_P3_RequestPending  0b1) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_READY_n  0b1)) (bv-comp P2_P1_P3_NA_n  0b0))   0b0)) ;5550
                                        if ((((P2_P1_P3_RequestPending == 1'b0) & (P2_P1_P3_HOLD == 1'b0)) & (P2_P1_P3_READY_n == 1'b0))) begin
                                            $display(";A 5552");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_RequestPending  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_READY_n  0b0))   0b1)) ;5552
                                            P2_P1_P3_State <= #1 3'sb001; $display(";A 5554");		//(= P2_P1_P3_State    0b001)) ;5554
                                        end
                                        else begin
                                            $display(";A 5553");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_RequestPending  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_READY_n  0b0))   0b0)) ;5553
                                            if (((P2_P1_P3_HOLD == 1'b1) & (P2_P1_P3_READY_n == 1'b1))) begin
                                                $display(";A 5555");		//(= (bv-and (bv-comp P2_P1_P3_HOLD  0b1) (bv-comp P2_P1_P3_READY_n  0b1))   0b1)) ;5555
                                                P2_P1_P3_State <= #1 3'sb101; $display(";A 5557");		//(= P2_P1_P3_State    0b101)) ;5557
                                            end
                                            else begin
                                                $display(";A 5556");		//(= (bv-and (bv-comp P2_P1_P3_HOLD  0b1) (bv-comp P2_P1_P3_READY_n  0b1))   0b0)) ;5556
                                                P2_P1_P3_State <= #1 3'sb011; $display(";A 5558");		//(= P2_P1_P3_State    0b011)) ;5558
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P2_P1_P3_StateBS16 <= #1 P2_P1_P3_BS16_n; $display(";A 5559");		//(= P2_P1_P3_StateBS16    P2_P1_P3_BS16_n )) ;5559
                        if ((P2_P1_P3_BS16_n == 1'b0)) begin
                            $display(";A 5560");		//(= (bv-comp P2_P1_P3_BS16_n  0b0)   0b1)) ;5560
                            P2_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 5562");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000001)) ;5562
                        end
                        else begin
                            $display(";A 5561");		//(= (bv-comp P2_P1_P3_BS16_n  0b0)   0b0)) ;5561
                            P2_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 5563");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;5563
                        end
                        P2_P1_P3_StateNA <= #1 P2_P1_P3_NA_n; $display(";A 5564");		//(= P2_P1_P3_StateNA    P2_P1_P3_NA_n )) ;5564
                        P2_P1_P3_ADS_n <= #1 1'b1; $display(";A 5565");		//(= P2_P1_P3_ADS_n    0b1)) ;5565
                    end
                3'b100 :
                    begin
                        $display(";A 5566");		//(= P2_P1_P3_State    0b100)) ;5566
                        if ((((P2_P1_P3_NA_n == 1'b0) & (P2_P1_P3_HOLD == 1'b0)) & (P2_P1_P3_RequestPending == 1'b1))) begin
                            $display(";A 5567");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_NA_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b1))   0b1)) ;5567
                            P2_P1_P3_State <= #1 3'sb110; $display(";A 5569");		//(= P2_P1_P3_State    0b110)) ;5569
                        end
                        else begin
                            $display(";A 5568");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_NA_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b1))   0b0)) ;5568
                            if (((P2_P1_P3_NA_n == 1'b0) & ((P2_P1_P3_HOLD == 1'b1) | (P2_P1_P3_RequestPending == 1'b0)))) begin
                                $display(";A 5570");		//(= (bv-and (bv-comp P2_P1_P3_NA_n  0b0) (bv-or (bv-comp P2_P1_P3_HOLD  0b1) (bv-comp P2_P1_P3_RequestPending  0b0)))   0b1)) ;5570
                                P2_P1_P3_State <= #1 3'sb111; $display(";A 5572");		//(= P2_P1_P3_State    0b111)) ;5572
                            end
                            else begin
                                $display(";A 5571");		//(= (bv-and (bv-comp P2_P1_P3_NA_n  0b0) (bv-or (bv-comp P2_P1_P3_HOLD  0b1) (bv-comp P2_P1_P3_RequestPending  0b0)))   0b0)) ;5571
                                if ((P2_P1_P3_NA_n == 1'b1)) begin
                                    $display(";A 5573");		//(= (bv-comp P2_P1_P3_NA_n  0b1)   0b1)) ;5573
                                    P2_P1_P3_State <= #1 3'sb011; $display(";A 5575");		//(= P2_P1_P3_State    0b011)) ;5575
                                end
                                else begin
                                    $display(";A 5574");		//(= (bv-comp P2_P1_P3_NA_n  0b1)   0b0)) ;5574
                                    P2_P1_P3_State <= #1 3'sb100; $display(";A 5576");		//(= P2_P1_P3_State    0b100)) ;5576
                                end
                            end
                        end
                        P2_P1_P3_StateBS16 <= #1 P2_P1_P3_BS16_n; $display(";A 5577");		//(= P2_P1_P3_StateBS16    P2_P1_P3_BS16_n )) ;5577
                        if ((P2_P1_P3_BS16_n == 1'b0)) begin
                            $display(";A 5578");		//(= (bv-comp P2_P1_P3_BS16_n  0b0)   0b1)) ;5578
                            P2_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 5580");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000001)) ;5580
                        end
                        else begin
                            $display(";A 5579");		//(= (bv-comp P2_P1_P3_BS16_n  0b0)   0b0)) ;5579
                            P2_P1_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 5581");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;5581
                        end
                        P2_P1_P3_StateNA <= #1 P2_P1_P3_NA_n; $display(";A 5582");		//(= P2_P1_P3_StateNA    P2_P1_P3_NA_n )) ;5582
                        P2_P1_P3_ADS_n <= #1 1'b1; $display(";A 5583");		//(= P2_P1_P3_ADS_n    0b1)) ;5583
                    end
                3'b101 :
                    begin
                        $display(";A 5584");		//(= P2_P1_P3_State    0b101)) ;5584
                        if (((P2_P1_P3_HOLD == 1'b0) & (P2_P1_P3_RequestPending == 1'b1))) begin
                            $display(";A 5585");		//(= (bv-and (bv-comp P2_P1_P3_HOLD  0b0) (bv-comp P2_P1_P3_RequestPending  0b1))   0b1)) ;5585
                            P2_P1_P3_State <= #1 3'sb010; $display(";A 5587");		//(= P2_P1_P3_State    0b010)) ;5587
                        end
                        else begin
                            $display(";A 5586");		//(= (bv-and (bv-comp P2_P1_P3_HOLD  0b0) (bv-comp P2_P1_P3_RequestPending  0b1))   0b0)) ;5586
                            if (((P2_P1_P3_HOLD == 1'b0) & (P2_P1_P3_RequestPending == 1'b0))) begin
                                $display(";A 5588");		//(= (bv-and (bv-comp P2_P1_P3_HOLD  0b0) (bv-comp P2_P1_P3_RequestPending  0b0))   0b1)) ;5588
                                P2_P1_P3_State <= #1 3'sb001; $display(";A 5590");		//(= P2_P1_P3_State    0b001)) ;5590
                            end
                            else begin
                                $display(";A 5589");		//(= (bv-and (bv-comp P2_P1_P3_HOLD  0b0) (bv-comp P2_P1_P3_RequestPending  0b0))   0b0)) ;5589
                                P2_P1_P3_State <= #1 3'sb101; $display(";A 5591");		//(= P2_P1_P3_State    0b101)) ;5591
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 5592");		//(= P2_P1_P3_State    0b110)) ;5592
                        P2_P1_P3_Address <= #1 ((P2_P1_P3_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 5593");		//(= P2_P1_P3_Address    (bv-smod (bv-sdiv P2_P1_P3_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;5593
                        P2_P1_P3_BE_n <= #1 P2_P1_P3_ByteEnable; $display(";A 5594");		//(= P2_P1_P3_BE_n    P2_P1_P3_ByteEnable )) ;5594
                        P2_P1_P3_M_IO_n <= #1 P2_P1_P3_MemoryFetch; $display(";A 5595");		//(= P2_P1_P3_M_IO_n    P2_P1_P3_MemoryFetch )) ;5595
                        if ((P2_P1_P3_ReadRequest == 1'b1)) begin
                            $display(";A 5596");		//(= (bv-comp P2_P1_P3_ReadRequest  0b1)   0b1)) ;5596
                            P2_P1_P3_W_R_n <= #1 1'b0; $display(";A 5598");		//(= P2_P1_P3_W_R_n    0b0)) ;5598
                        end
                        else begin
                            $display(";A 5597");		//(= (bv-comp P2_P1_P3_ReadRequest  0b1)   0b0)) ;5597
                            P2_P1_P3_W_R_n <= #1 1'b1; $display(";A 5599");		//(= P2_P1_P3_W_R_n    0b1)) ;5599
                        end
                        if ((P2_P1_P3_CodeFetch == 1'b1)) begin
                            $display(";A 5600");		//(= (bv-comp P2_P1_P3_CodeFetch  0b1)   0b1)) ;5600
                            P2_P1_P3_D_C_n <= #1 1'b0; $display(";A 5602");		//(= P2_P1_P3_D_C_n    0b0)) ;5602
                        end
                        else begin
                            $display(";A 5601");		//(= (bv-comp P2_P1_P3_CodeFetch  0b1)   0b0)) ;5601
                            P2_P1_P3_D_C_n <= #1 1'b1; $display(";A 5603");		//(= P2_P1_P3_D_C_n    0b1)) ;5603
                        end
                        P2_P1_P3_ADS_n <= #1 1'b0; $display(";A 5604");		//(= P2_P1_P3_ADS_n    0b0)) ;5604
                        if ((P2_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 5605");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5605
                            P2_P1_P3_State <= #1 3'sb100; $display(";A 5607");		//(= P2_P1_P3_State    0b100)) ;5607
                        end
                        else begin
                            $display(";A 5606");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5606
                            P2_P1_P3_State <= #1 3'sb110; $display(";A 5608");		//(= P2_P1_P3_State    0b110)) ;5608
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 5609");		//(= P2_P1_P3_State    0b111)) ;5609
                        if ((((P2_P1_P3_READY_n == 1'b1) & (P2_P1_P3_RequestPending == 1'b1)) & (P2_P1_P3_HOLD == 1'b0))) begin
                            $display(";A 5610");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b1) (bv-comp P2_P1_P3_RequestPending  0b1)) (bv-comp P2_P1_P3_HOLD  0b0))   0b1)) ;5610
                            P2_P1_P3_State <= #1 3'sb110; $display(";A 5612");		//(= P2_P1_P3_State    0b110)) ;5612
                        end
                        else begin
                            $display(";A 5611");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b1) (bv-comp P2_P1_P3_RequestPending  0b1)) (bv-comp P2_P1_P3_HOLD  0b0))   0b0)) ;5611
                            if (((P2_P1_P3_READY_n == 1'b0) & (P2_P1_P3_HOLD == 1'b1))) begin
                                $display(";A 5613");		//(= (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b1))   0b1)) ;5613
                                P2_P1_P3_State <= #1 3'sb101; $display(";A 5615");		//(= P2_P1_P3_State    0b101)) ;5615
                            end
                            else begin
                                $display(";A 5614");		//(= (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b1))   0b0)) ;5614
                                if ((((P2_P1_P3_READY_n == 1'b0) & (P2_P1_P3_HOLD == 1'b0)) & (P2_P1_P3_RequestPending == 1'b1))) begin
                                    $display(";A 5616");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b1))   0b1)) ;5616
                                    P2_P1_P3_State <= #1 3'sb010; $display(";A 5618");		//(= P2_P1_P3_State    0b010)) ;5618
                                end
                                else begin
                                    $display(";A 5617");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b1))   0b0)) ;5617
                                    if ((((P2_P1_P3_READY_n == 1'b0) & (P2_P1_P3_HOLD == 1'b0)) & (P2_P1_P3_RequestPending == 1'b0))) begin
                                        $display(";A 5619");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b0))   0b1)) ;5619
                                        P2_P1_P3_State <= #1 3'sb001; $display(";A 5621");		//(= P2_P1_P3_State    0b001)) ;5621
                                    end
                                    else begin
                                        $display(";A 5620");		//(= (bv-and (bv-and (bv-comp P2_P1_P3_READY_n  0b0) (bv-comp P2_P1_P3_HOLD  0b0)) (bv-comp P2_P1_P3_RequestPending  0b0))   0b0)) ;5620
                                        P2_P1_P3_State <= #1 3'sb111; $display(";A 5622");		//(= P2_P1_P3_State    0b111)) ;5622
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:8577
    always @(posedge P2_P1_P3_RESET or posedge P2_P1_P3_CLOCK) begin
        if ((P2_P1_P3_RESET == 1'b1)) begin
            $display(";A 5623");		//(= (bv-comp P2_P1_P3_RESET  0b1)   0b1)) ;5623
            P2_P1_P3_State2 = 4'sb0000; $display(";A 5625");		//(= P2_P1_P3_State2    0b0000)) ;5625
            P2_P1_P3_InstQueue[0] = 8'b00000000; $display(";A 5626");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5626
            P2_P1_P3_InstQueue[1] = 8'b00000000; $display(";A 5627");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5627
            P2_P1_P3_InstQueue[2] = 8'b00000000; $display(";A 5628");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5628
            P2_P1_P3_InstQueue[3] = 8'b00000000; $display(";A 5629");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5629
            P2_P1_P3_InstQueue[4] = 8'b00000000; $display(";A 5630");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5630
            P2_P1_P3_InstQueue[5] = 8'b00000000; $display(";A 5631");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5631
            P2_P1_P3_InstQueue[6] = 8'b00000000; $display(";A 5632");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5632
            P2_P1_P3_InstQueue[7] = 8'b00000000; $display(";A 5633");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5633
            P2_P1_P3_InstQueue[8] = 8'b00000000; $display(";A 5634");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5634
            P2_P1_P3_InstQueue[9] = 8'b00000000; $display(";A 5635");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5635
            P2_P1_P3_InstQueue[10] = 8'b00000000; $display(";A 5636");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5636
            P2_P1_P3_InstQueue[11] = 8'b00000000; $display(";A 5637");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5637
            P2_P1_P3_InstQueue[12] = 8'b00000000; $display(";A 5638");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5638
            P2_P1_P3_InstQueue[13] = 8'b00000000; $display(";A 5639");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5639
            P2_P1_P3_InstQueue[14] = 8'b00000000; $display(";A 5640");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5640
            P2_P1_P3_InstQueue[15] = 8'b00000000; $display(";A 5641");		//(= P2_P1_P3_InstQueue    0b00000000)) ;5641
            P2_P1_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 5642");		//(= P2_P1_P3_InstQueueRd_Addr    0b00000)) ;5642
            P2_P1_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 5643");		//(= P2_P1_P3_InstQueueWr_Addr    0b00000)) ;5643
            P2_P1_P3_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 5644");		//(= P2_P1_P3_InstAddrPointer    0b00000000000000000000000000000000)) ;5644
            P2_P1_P3_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 5645");		//(= P2_P1_P3_PhyAddrPointer    0b00000000000000000000000000000000)) ;5645
            P2_P1_P3_Extended = 1'b0; $display(";A 5646");		//(= P2_P1_P3_Extended    0b0)) ;5646
            P2_P1_P3_More = 1'b0; $display(";A 5647");		//(= P2_P1_P3_More    0b0)) ;5647
            P2_P1_P3_Flush = 1'b0; $display(";A 5648");		//(= P2_P1_P3_Flush    0b0)) ;5648
            P2_P1_P3_lWord = 16'sb0000000000000000; $display(";A 5649");		//(= P2_P1_P3_lWord    0b0000000000000000)) ;5649
            P2_P1_P3_uWord = 15'sb000000000000000; $display(";A 5650");		//(= P2_P1_P3_uWord    0b000000000000000)) ;5650
            P2_P1_P3_fWord = 32'sb00000000000000000000000000000000; $display(";A 5651");		//(= P2_P1_P3_fWord    0b00000000000000000000000000000000)) ;5651
            P2_P1_P3_CodeFetch <= #1 1'b0; $display(";A 5652");		//(= P2_P1_P3_CodeFetch    0b0)) ;5652
            P2_P1_P3_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 5653");		//(= P2_P1_P3_Datao    0b00000000000000000000000000000000)) ;5653
            P2_P1_P3_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 5654");		//(= P2_P1_P3_EAX    0b00000000000000000000000000000000)) ;5654
            P2_P1_P3_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 5655");		//(= P2_P1_P3_EBX    0b00000000000000000000000000000000)) ;5655
            P2_P1_P3_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 5656");		//(= P2_P1_P3_rEIP    0b00000000000000000000000000000000)) ;5656
            P2_P1_P3_ReadRequest <= #1 1'b0; $display(";A 5657");		//(= P2_P1_P3_ReadRequest    0b0)) ;5657
            P2_P1_P3_MemoryFetch <= #1 1'b0; $display(";A 5658");		//(= P2_P1_P3_MemoryFetch    0b0)) ;5658
            P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5659");		//(= P2_P1_P3_RequestPending    0b0)) ;5659
        end
        else begin
            $display(";A 5624");		//(= (bv-comp P2_P1_P3_RESET  0b1)   0b0)) ;5624
            case (P2_P1_P3_State2)
                4'b0000 :
                    begin
                        $display(";A 5660");		//(= P2_P1_P3_State2    0b0000)) ;5660
                        P2_P1_P3_PhyAddrPointer = P2_P1_P3_rEIP; $display(";A 5661");		//(= P2_P1_P3_PhyAddrPointer    P2_P1_P3_rEIP )) ;5661
                        P2_P1_P3_InstAddrPointer = P2_P1_P3_PhyAddrPointer; $display(";A 5662");		//(= P2_P1_P3_InstAddrPointer    P2_P1_P3_PhyAddrPointer )) ;5662
                        P2_P1_P3_State2 = 4'sb0001; $display(";A 5663");		//(= P2_P1_P3_State2    0b0001)) ;5663
                        P2_P1_P3_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 5664");		//(= P2_P1_P3_rEIP    0b00000000000011111111111111110000)) ;5664
                        P2_P1_P3_ReadRequest <= #1 1'b1; $display(";A 5665");		//(= P2_P1_P3_ReadRequest    0b1)) ;5665
                        P2_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 5666");		//(= P2_P1_P3_MemoryFetch    0b1)) ;5666
                        P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5667");		//(= P2_P1_P3_RequestPending    0b1)) ;5667
                    end
                4'b0001 :
                    begin
                        $display(";A 5668");		//(= P2_P1_P3_State2    0b0001)) ;5668
                        P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5669");		//(= P2_P1_P3_RequestPending    0b1)) ;5669
                        P2_P1_P3_ReadRequest <= #1 1'b1; $display(";A 5670");		//(= P2_P1_P3_ReadRequest    0b1)) ;5670
                        P2_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 5671");		//(= P2_P1_P3_MemoryFetch    0b1)) ;5671
                        P2_P1_P3_CodeFetch <= #1 1'b1; $display(";A 5672");		//(= P2_P1_P3_CodeFetch    0b1)) ;5672
                        if ((P2_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 5673");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5673
                            P2_P1_P3_State2 = 4'sb0010; $display(";A 5675");		//(= P2_P1_P3_State2    0b0010)) ;5675
                        end
                        else begin
                            $display(";A 5674");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5674
                            P2_P1_P3_State2 = 4'sb0001; $display(";A 5676");		//(= P2_P1_P3_State2    0b0001)) ;5676
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 5677");		//(= P2_P1_P3_State2    0b0010)) ;5677
                        P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5678");		//(= P2_P1_P3_RequestPending    0b0)) ;5678
                        P2_P1_P3_InstQueue[P2_P1_P3_InstQueueWr_Addr] = (P2_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 5679");		//(= P2_P1_P3_InstQueue    (bv-smod P2_P1_P3_Datai  0b00000000000000000000000100000000))) ;5679
                        P2_P1_P3_InstQueueWr_Addr = ((P2_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5680");		//(= P2_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5680
                        P2_P1_P3_InstQueue[P2_P1_P3_InstQueueWr_Addr] = (P2_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 5681");		//(= P2_P1_P3_InstQueue    (bv-smod P2_P1_P3_Datai  0b00000000000000000000000100000000))) ;5681
                        P2_P1_P3_InstQueueWr_Addr = ((P2_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5682");		//(= P2_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5682
                        if ((P2_P1_P3_StateBS16 == 1'b1)) begin
                            $display(";A 5683");		//(= (bv-comp P2_P1_P3_StateBS16  0b1)   0b1)) ;5683
                            P2_P1_P3_InstQueue[P2_P1_P3_InstQueueWr_Addr] = ((P2_P1_P3_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 5685");		//(= P2_P1_P3_InstQueue    (bv-smod (bv-sdiv P2_P1_P3_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;5685
                            P2_P1_P3_InstQueueWr_Addr = ((P2_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5686");		//(= P2_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5686
                            P2_P1_P3_InstQueue[P2_P1_P3_InstQueueWr_Addr] = ((P2_P1_P3_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 5687");		//(= P2_P1_P3_InstQueue    (bv-smod (bv-sdiv P2_P1_P3_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;5687
                            P2_P1_P3_InstQueueWr_Addr = ((P2_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5688");		//(= P2_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5688
                            P2_P1_P3_PhyAddrPointer = (P2_P1_P3_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 5689");		//(= P2_P1_P3_PhyAddrPointer    (bv-add P2_P1_P3_PhyAddrPointer  0b00000000000000000000000000000100))) ;5689
                            P2_P1_P3_State2 = 4'sb0101; $display(";A 5690");		//(= P2_P1_P3_State2    0b0101)) ;5690
                        end
                        else begin
                            $display(";A 5684");		//(= (bv-comp P2_P1_P3_StateBS16  0b1)   0b0)) ;5684
                            P2_P1_P3_PhyAddrPointer = (P2_P1_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5691");		//(= P2_P1_P3_PhyAddrPointer    (bv-add P2_P1_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;5691
                            if ((P2_P1_P3_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 5692");		//(= (bool-to-bv (bv-slt P2_P1_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;5692
                                P2_P1_P3_rEIP <= #1 (-P2_P1_P3_PhyAddrPointer); $display(";A 5694");		//(= P2_P1_P3_rEIP    (bv-neg P2_P1_P3_PhyAddrPointer ))) ;5694
                            end
                            else begin
                                $display(";A 5693");		//(= (bool-to-bv (bv-slt P2_P1_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;5693
                                P2_P1_P3_rEIP <= #1 P2_P1_P3_PhyAddrPointer; $display(";A 5695");		//(= P2_P1_P3_rEIP    P2_P1_P3_PhyAddrPointer )) ;5695
                            end
                            P2_P1_P3_State2 = 4'sb0011; $display(";A 5696");		//(= P2_P1_P3_State2    0b0011)) ;5696
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 5697");		//(= P2_P1_P3_State2    0b0011)) ;5697
                        P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5698");		//(= P2_P1_P3_RequestPending    0b1)) ;5698
                        if ((P2_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 5699");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5699
                            P2_P1_P3_State2 = 4'sb0100; $display(";A 5701");		//(= P2_P1_P3_State2    0b0100)) ;5701
                        end
                        else begin
                            $display(";A 5700");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5700
                            P2_P1_P3_State2 = 4'sb0011; $display(";A 5702");		//(= P2_P1_P3_State2    0b0011)) ;5702
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 5703");		//(= P2_P1_P3_State2    0b0100)) ;5703
                        P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5704");		//(= P2_P1_P3_RequestPending    0b0)) ;5704
                        P2_P1_P3_InstQueue[P2_P1_P3_InstQueueWr_Addr] = (P2_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 5705");		//(= P2_P1_P3_InstQueue    (bv-smod P2_P1_P3_Datai  0b00000000000000000000000100000000))) ;5705
                        P2_P1_P3_InstQueueWr_Addr = ((P2_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5706");		//(= P2_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5706
                        P2_P1_P3_InstQueue[P2_P1_P3_InstQueueWr_Addr] = (P2_P1_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 5707");		//(= P2_P1_P3_InstQueue    (bv-smod P2_P1_P3_Datai  0b00000000000000000000000100000000))) ;5707
                        P2_P1_P3_InstQueueWr_Addr = ((P2_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5708");		//(= P2_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5708
                        P2_P1_P3_PhyAddrPointer = (P2_P1_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5709");		//(= P2_P1_P3_PhyAddrPointer    (bv-add P2_P1_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;5709
                        P2_P1_P3_State2 = 4'sb0101; $display(";A 5710");		//(= P2_P1_P3_State2    0b0101)) ;5710
                    end
                4'b0101 :
                    begin
                        $display(";A 5711");		//(= P2_P1_P3_State2    0b0101)) ;5711
                        case (P2_P1_P3_InstQueue[P2_P1_P3_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 5712");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b10010000)) ;5712
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5713");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5713
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5714");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5714
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5715");		//(= P2_P1_P3_Flush    0b0)) ;5715
                                    P2_P1_P3_More = 1'b0; $display(";A 5716");		//(= P2_P1_P3_More    0b0)) ;5716
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 5717");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b01100110)) ;5717
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5718");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5718
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5719");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5719
                                    P2_P1_P3_Extended = 1'b1; $display(";A 5720");		//(= P2_P1_P3_Extended    0b1)) ;5720
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5721");		//(= P2_P1_P3_Flush    0b0)) ;5721
                                    P2_P1_P3_More = 1'b0; $display(";A 5722");		//(= P2_P1_P3_More    0b0)) ;5722
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 5723");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b11101011)) ;5723
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 5724");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;5724
                                        if ((P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 5726");		//(= (bool-to-bv (bv-gt P2_P1_P3_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;5726
                                            P2_P1_P3_PhyAddrPointer = ((P2_P1_P3_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 5728");		//(= P2_P1_P3_PhyAddrPointer    (bv-sub (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P2_P1_P3_InstQueue 0 )))) ;5728
                                            P2_P1_P3_InstAddrPointer = P2_P1_P3_PhyAddrPointer; $display(";A 5729");		//(= P2_P1_P3_InstAddrPointer    P2_P1_P3_PhyAddrPointer )) ;5729
                                        end
                                        else begin
                                            $display(";A 5727");		//(= (bool-to-bv (bv-gt P2_P1_P3_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;5727
                                            P2_P1_P3_PhyAddrPointer = ((P2_P1_P3_InstAddrPointer + 32'b00000000000000000000000000000010) + P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 5730");		//(= P2_P1_P3_PhyAddrPointer    (bv-add (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000010) P2_P1_P3_InstQueue 0 ))) ;5730
                                            P2_P1_P3_InstAddrPointer = P2_P1_P3_PhyAddrPointer; $display(";A 5731");		//(= P2_P1_P3_InstAddrPointer    P2_P1_P3_PhyAddrPointer )) ;5731
                                        end
                                        P2_P1_P3_Flush = 1'b1; $display(";A 5732");		//(= P2_P1_P3_Flush    0b1)) ;5732
                                        P2_P1_P3_More = 1'b0; $display(";A 5733");		//(= P2_P1_P3_More    0b0)) ;5733
                                    end
                                    else begin
                                        $display(";A 5725");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;5725
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5734");		//(= P2_P1_P3_Flush    0b0)) ;5734
                                        P2_P1_P3_More = 1'b1; $display(";A 5735");		//(= P2_P1_P3_More    0b1)) ;5735
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 5736");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b11101001)) ;5736
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 5737");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;5737
                                        P2_P1_P3_PhyAddrPointer = ((P2_P1_P3_InstAddrPointer + 32'b00000000000000000000000000000101) + P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 5739");		//(= P2_P1_P3_PhyAddrPointer    (bv-add (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000101) P2_P1_P3_InstQueue 0 ))) ;5739
                                        P2_P1_P3_InstAddrPointer = P2_P1_P3_PhyAddrPointer; $display(";A 5740");		//(= P2_P1_P3_InstAddrPointer    P2_P1_P3_PhyAddrPointer )) ;5740
                                        P2_P1_P3_Flush = 1'b1; $display(";A 5741");		//(= P2_P1_P3_Flush    0b1)) ;5741
                                        P2_P1_P3_More = 1'b0; $display(";A 5742");		//(= P2_P1_P3_More    0b0)) ;5742
                                    end
                                    else begin
                                        $display(";A 5738");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;5738
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5743");		//(= P2_P1_P3_Flush    0b0)) ;5743
                                        P2_P1_P3_More = 1'b1; $display(";A 5744");		//(= P2_P1_P3_More    0b1)) ;5744
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 5745");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b11101010)) ;5745
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5746");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5746
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5747");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5747
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5748");		//(= P2_P1_P3_Flush    0b0)) ;5748
                                    P2_P1_P3_More = 1'b0; $display(";A 5749");		//(= P2_P1_P3_More    0b0)) ;5749
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 5750");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b10110000)) ;5750
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5751");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5751
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5752");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5752
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5753");		//(= P2_P1_P3_Flush    0b0)) ;5753
                                    P2_P1_P3_More = 1'b0; $display(";A 5754");		//(= P2_P1_P3_More    0b0)) ;5754
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 5755");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b10111000)) ;5755
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 5756");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;5756
                                        P2_P1_P3_EAX <= #1 ((((P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 5758");		//(= P2_P1_P3_EAX    (bv-add (bv-add (bv-add (bv-mul P2_P1_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P1_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P1_P3_InstQueue 0  0b00000000000000000000000100000000)) P2_P1_P3_InstQueue 0 ))) ;5758
                                        P2_P1_P3_More = 1'b0; $display(";A 5759");		//(= P2_P1_P3_More    0b0)) ;5759
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5760");		//(= P2_P1_P3_Flush    0b0)) ;5760
                                        P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 5761");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;5761
                                        P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 5762");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;5762
                                    end
                                    else begin
                                        $display(";A 5757");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;5757
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5763");		//(= P2_P1_P3_Flush    0b0)) ;5763
                                        P2_P1_P3_More = 1'b1; $display(";A 5764");		//(= P2_P1_P3_More    0b1)) ;5764
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 5765");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b10111011)) ;5765
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 5766");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;5766
                                        P2_P1_P3_EBX <= #1 ((((P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P1_P3_InstQueue[((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 5768");		//(= P2_P1_P3_EBX    (bv-add (bv-add (bv-add (bv-mul P2_P1_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P1_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P1_P3_InstQueue 0  0b00000000000000000000000100000000)) P2_P1_P3_InstQueue 0 ))) ;5768
                                        P2_P1_P3_More = 1'b0; $display(";A 5769");		//(= P2_P1_P3_More    0b0)) ;5769
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5770");		//(= P2_P1_P3_Flush    0b0)) ;5770
                                        P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 5771");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;5771
                                        P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 5772");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;5772
                                    end
                                    else begin
                                        $display(";A 5767");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;5767
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5773");		//(= P2_P1_P3_Flush    0b0)) ;5773
                                        P2_P1_P3_More = 1'b1; $display(";A 5774");		//(= P2_P1_P3_More    0b1)) ;5774
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 5775");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b10001011)) ;5775
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5776");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5776
                                        if ((P2_P1_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 5778");		//(= (bool-to-bv (bv-slt P2_P1_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;5778
                                            P2_P1_P3_rEIP <= #1 (-P2_P1_P3_EBX); $display(";A 5780");		//(= P2_P1_P3_rEIP    (bv-neg P2_P1_P3_EBX ))) ;5780
                                        end
                                        else begin
                                            $display(";A 5779");		//(= (bool-to-bv (bv-slt P2_P1_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;5779
                                            P2_P1_P3_rEIP <= #1 P2_P1_P3_EBX; $display(";A 5781");		//(= P2_P1_P3_rEIP    P2_P1_P3_EBX )) ;5781
                                        end
                                        P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5782");		//(= P2_P1_P3_RequestPending    0b1)) ;5782
                                        P2_P1_P3_ReadRequest <= #1 1'b1; $display(";A 5783");		//(= P2_P1_P3_ReadRequest    0b1)) ;5783
                                        P2_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 5784");		//(= P2_P1_P3_MemoryFetch    0b1)) ;5784
                                        P2_P1_P3_CodeFetch <= #1 1'b0; $display(";A 5785");		//(= P2_P1_P3_CodeFetch    0b0)) ;5785
                                        if ((P2_P1_P3_READY_n == 1'b0)) begin
                                            $display(";A 5786");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5786
                                            P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5788");		//(= P2_P1_P3_RequestPending    0b0)) ;5788
                                            P2_P1_P3_uWord = (P2_P1_P3_Datai % 32'b00000000000000001000000000000000); $display(";A 5789");		//(= P2_P1_P3_uWord    (bv-smod P2_P1_P3_Datai  0b00000000000000001000000000000000))) ;5789
                                            if ((P2_P1_P3_StateBS16 == 1'b1)) begin
                                                $display(";A 5790");		//(= (bv-comp P2_P1_P3_StateBS16  0b1)   0b1)) ;5790
                                                P2_P1_P3_lWord = (P2_P1_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 5792");		//(= P2_P1_P3_lWord    (bv-smod P2_P1_P3_Datai  0b00000000000000010000000000000000))) ;5792
                                            end
                                            else begin
                                                $display(";A 5791");		//(= (bv-comp P2_P1_P3_StateBS16  0b1)   0b0)) ;5791
                                                P2_P1_P3_rEIP <= #1 (P2_P1_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 5793");		//(= P2_P1_P3_rEIP    (bv-add P2_P1_P3_rEIP  0b00000000000000000000000000000010))) ;5793
                                                P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5794");		//(= P2_P1_P3_RequestPending    0b1)) ;5794
                                                if ((P2_P1_P3_READY_n == 1'b0)) begin
                                                    $display(";A 5795");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5795
                                                    P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5797");		//(= P2_P1_P3_RequestPending    0b0)) ;5797
                                                    P2_P1_P3_lWord = (P2_P1_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 5798");		//(= P2_P1_P3_lWord    (bv-smod P2_P1_P3_Datai  0b00000000000000010000000000000000))) ;5798
                                                end
                                                else begin
                                                    $display(";A 5796");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5796
                                                end
                                            end
                                            if ((P2_P1_P3_READY_n == 1'b0)) begin
                                                $display(";A 5799");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5799
                                                P2_P1_P3_EAX <= #1 ((P2_P1_P3_uWord * 32'b00000000000000010000000000000000) + P2_P1_P3_lWord); $display(";A 5801");		//(= P2_P1_P3_EAX    (bv-add (bv-mul P2_P1_P3_uWord  0b00000000000000010000000000000000) P2_P1_P3_lWord ))) ;5801
                                                P2_P1_P3_More = 1'b0; $display(";A 5802");		//(= P2_P1_P3_More    0b0)) ;5802
                                                P2_P1_P3_Flush = 1'b0; $display(";A 5803");		//(= P2_P1_P3_Flush    0b0)) ;5803
                                                P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5804");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;5804
                                                P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5805");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5805
                                            end
                                            else begin
                                                $display(";A 5800");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5800
                                            end
                                        end
                                        else begin
                                            $display(";A 5787");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5787
                                        end
                                    end
                                    else begin
                                        $display(";A 5777");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5777
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5806");		//(= P2_P1_P3_Flush    0b0)) ;5806
                                        P2_P1_P3_More = 1'b1; $display(";A 5807");		//(= P2_P1_P3_More    0b1)) ;5807
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 5808");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b10001001)) ;5808
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5809");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5809
                                        if ((P2_P1_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 5811");		//(= (bool-to-bv (bv-slt P2_P1_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;5811
                                            P2_P1_P3_rEIP <= #1 P2_P1_P3_EBX; $display(";A 5813");		//(= P2_P1_P3_rEIP    P2_P1_P3_EBX )) ;5813
                                        end
                                        else begin
                                            $display(";A 5812");		//(= (bool-to-bv (bv-slt P2_P1_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;5812
                                            P2_P1_P3_rEIP <= #1 P2_P1_P3_EBX; $display(";A 5814");		//(= P2_P1_P3_rEIP    P2_P1_P3_EBX )) ;5814
                                        end
                                        P2_P1_P3_lWord = (P2_P1_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 5815");		//(= P2_P1_P3_lWord    (bv-smod P2_P1_P3_EAX  0b00000000000000010000000000000000))) ;5815
                                        P2_P1_P3_uWord = ((P2_P1_P3_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 5816");		//(= P2_P1_P3_uWord    (bv-smod (bv-sdiv P2_P1_P3_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;5816
                                        P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5817");		//(= P2_P1_P3_RequestPending    0b1)) ;5817
                                        P2_P1_P3_ReadRequest <= #1 1'b0; $display(";A 5818");		//(= P2_P1_P3_ReadRequest    0b0)) ;5818
                                        P2_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 5819");		//(= P2_P1_P3_MemoryFetch    0b1)) ;5819
                                        P2_P1_P3_CodeFetch <= #1 1'b0; $display(";A 5820");		//(= P2_P1_P3_CodeFetch    0b0)) ;5820
                                        if (((P2_P1_P3_State == 32'b00000000000000000000000000000010) | (P2_P1_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 5821");		//(= (bv-or (bv-comp P2_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P3_State  0b00000000000000000000000000000100))   0b1)) ;5821
                                            P2_P1_P3_Datao <= #1 ((P2_P1_P3_uWord * 32'b00000000000000010000000000000000) + P2_P1_P3_lWord); $display(";A 5823");		//(= P2_P1_P3_Datao    (bv-add (bv-mul P2_P1_P3_uWord  0b00000000000000010000000000000000) P2_P1_P3_lWord ))) ;5823
                                            if ((P2_P1_P3_READY_n == 1'b0)) begin
                                                $display(";A 5824");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5824
                                                P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5826");		//(= P2_P1_P3_RequestPending    0b0)) ;5826
                                                if ((P2_P1_P3_StateBS16 == 1'b0)) begin
                                                    $display(";A 5827");		//(= (bv-comp P2_P1_P3_StateBS16  0b0)   0b1)) ;5827
                                                    P2_P1_P3_rEIP <= #1 (P2_P1_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 5829");		//(= P2_P1_P3_rEIP    (bv-add P2_P1_P3_rEIP  0b00000000000000000000000000000010))) ;5829
                                                    P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5830");		//(= P2_P1_P3_RequestPending    0b1)) ;5830
                                                    P2_P1_P3_ReadRequest <= #1 1'b0; $display(";A 5831");		//(= P2_P1_P3_ReadRequest    0b0)) ;5831
                                                    P2_P1_P3_MemoryFetch <= #1 1'b1; $display(";A 5832");		//(= P2_P1_P3_MemoryFetch    0b1)) ;5832
                                                    P2_P1_P3_CodeFetch <= #1 1'b0; $display(";A 5833");		//(= P2_P1_P3_CodeFetch    0b0)) ;5833
                                                    P2_P1_P3_State2 = 4'sb0110; $display(";A 5834");		//(= P2_P1_P3_State2    0b0110)) ;5834
                                                end
                                                else begin
                                                    $display(";A 5828");		//(= (bv-comp P2_P1_P3_StateBS16  0b0)   0b0)) ;5828
                                                end
                                                P2_P1_P3_More = 1'b0; $display(";A 5835");		//(= P2_P1_P3_More    0b0)) ;5835
                                                P2_P1_P3_Flush = 1'b0; $display(";A 5836");		//(= P2_P1_P3_Flush    0b0)) ;5836
                                                P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5837");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;5837
                                                P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5838");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5838
                                            end
                                            else begin
                                                $display(";A 5825");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5825
                                            end
                                        end
                                        else begin
                                            $display(";A 5822");		//(= (bv-or (bv-comp P2_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P3_State  0b00000000000000000000000000000100))   0b0)) ;5822
                                        end
                                    end
                                    else begin
                                        $display(";A 5810");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5810
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5839");		//(= P2_P1_P3_Flush    0b0)) ;5839
                                        P2_P1_P3_More = 1'b1; $display(";A 5840");		//(= P2_P1_P3_More    0b1)) ;5840
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 5841");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b11100100)) ;5841
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5842");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5842
                                        P2_P1_P3_rEIP <= #1 (P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 5844");		//(= P2_P1_P3_rEIP    (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;5844
                                        P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5845");		//(= P2_P1_P3_RequestPending    0b1)) ;5845
                                        P2_P1_P3_ReadRequest <= #1 1'b1; $display(";A 5846");		//(= P2_P1_P3_ReadRequest    0b1)) ;5846
                                        P2_P1_P3_MemoryFetch <= #1 1'b0; $display(";A 5847");		//(= P2_P1_P3_MemoryFetch    0b0)) ;5847
                                        P2_P1_P3_CodeFetch <= #1 1'b0; $display(";A 5848");		//(= P2_P1_P3_CodeFetch    0b0)) ;5848
                                        if ((P2_P1_P3_READY_n == 1'b0)) begin
                                            $display(";A 5849");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5849
                                            P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5851");		//(= P2_P1_P3_RequestPending    0b0)) ;5851
                                            P2_P1_P3_EAX <= #1 P2_P1_P3_Datai; $display(";A 5852");		//(= P2_P1_P3_EAX    P2_P1_P3_Datai )) ;5852
                                            P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5853");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;5853
                                            P2_P1_P3_InstQueueRd_Addr = (P2_P1_P3_InstQueueRd_Addr + 5'b00010); $display(";A 5854");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-add P2_P1_P3_InstQueueRd_Addr  0b00010))) ;5854
                                            P2_P1_P3_Flush = 1'b0; $display(";A 5855");		//(= P2_P1_P3_Flush    0b0)) ;5855
                                            P2_P1_P3_More = 1'b0; $display(";A 5856");		//(= P2_P1_P3_More    0b0)) ;5856
                                        end
                                        else begin
                                            $display(";A 5850");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5850
                                        end
                                    end
                                    else begin
                                        $display(";A 5843");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5843
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5857");		//(= P2_P1_P3_Flush    0b0)) ;5857
                                        P2_P1_P3_More = 1'b1; $display(";A 5858");		//(= P2_P1_P3_More    0b1)) ;5858
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 5859");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b11100110)) ;5859
                                    if (((P2_P1_P3_InstQueueWr_Addr - P2_P1_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 5860");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;5860
                                        P2_P1_P3_rEIP <= #1 (P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 5862");		//(= P2_P1_P3_rEIP    (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;5862
                                        P2_P1_P3_RequestPending <= #1 1'b1; $display(";A 5863");		//(= P2_P1_P3_RequestPending    0b1)) ;5863
                                        P2_P1_P3_ReadRequest <= #1 1'b0; $display(";A 5864");		//(= P2_P1_P3_ReadRequest    0b0)) ;5864
                                        P2_P1_P3_MemoryFetch <= #1 1'b0; $display(";A 5865");		//(= P2_P1_P3_MemoryFetch    0b0)) ;5865
                                        P2_P1_P3_CodeFetch <= #1 1'b0; $display(";A 5866");		//(= P2_P1_P3_CodeFetch    0b0)) ;5866
                                        if (((P2_P1_P3_State == 32'b00000000000000000000000000000010) | (P2_P1_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 5867");		//(= (bv-or (bv-comp P2_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P3_State  0b00000000000000000000000000000100))   0b1)) ;5867
                                            P2_P1_P3_fWord = (P2_P1_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 5869");		//(= P2_P1_P3_fWord    (bv-smod P2_P1_P3_EAX  0b00000000000000010000000000000000))) ;5869
                                            P2_P1_P3_Datao <= #1 P2_P1_P3_fWord; $display(";A 5870");		//(= P2_P1_P3_Datao    P2_P1_P3_fWord )) ;5870
                                            if ((P2_P1_P3_READY_n == 1'b0)) begin
                                                $display(";A 5871");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5871
                                                P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5873");		//(= P2_P1_P3_RequestPending    0b0)) ;5873
                                                P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5874");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;5874
                                                P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5875");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5875
                                                P2_P1_P3_Flush = 1'b0; $display(";A 5876");		//(= P2_P1_P3_Flush    0b0)) ;5876
                                                P2_P1_P3_More = 1'b0; $display(";A 5877");		//(= P2_P1_P3_More    0b0)) ;5877
                                            end
                                            else begin
                                                $display(";A 5872");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5872
                                            end
                                        end
                                        else begin
                                            $display(";A 5868");		//(= (bv-or (bv-comp P2_P1_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P1_P3_State  0b00000000000000000000000000000100))   0b0)) ;5868
                                        end
                                    end
                                    else begin
                                        $display(";A 5861");		//(= (bool-to-bv (bv-ge (bv-sub P2_P1_P3_InstQueueWr_Addr  P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;5861
                                        P2_P1_P3_Flush = 1'b0; $display(";A 5878");		//(= P2_P1_P3_Flush    0b0)) ;5878
                                        P2_P1_P3_More = 1'b1; $display(";A 5879");		//(= P2_P1_P3_More    0b1)) ;5879
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 5880");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b00000100)) ;5880
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5881");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5881
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5882");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5882
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5883");		//(= P2_P1_P3_Flush    0b0)) ;5883
                                    P2_P1_P3_More = 1'b0; $display(";A 5884");		//(= P2_P1_P3_More    0b0)) ;5884
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 5885");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b00000101)) ;5885
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5886");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5886
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5887");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5887
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5888");		//(= P2_P1_P3_Flush    0b0)) ;5888
                                    P2_P1_P3_More = 1'b0; $display(";A 5889");		//(= P2_P1_P3_More    0b0)) ;5889
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 5890");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b11010000)) ;5890
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5891");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;5891
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5892");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5892
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5893");		//(= P2_P1_P3_Flush    0b0)) ;5893
                                    P2_P1_P3_More = 1'b0; $display(";A 5894");		//(= P2_P1_P3_More    0b0)) ;5894
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 5895");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b11000000)) ;5895
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 5896");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;5896
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 5897");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;5897
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5898");		//(= P2_P1_P3_Flush    0b0)) ;5898
                                    P2_P1_P3_More = 1'b0; $display(";A 5899");		//(= P2_P1_P3_More    0b0)) ;5899
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 5900");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b01000000)) ;5900
                                    P2_P1_P3_EAX <= #1 (P2_P1_P3_EAX + 32'sb00000000000000000000000000000001); $display(";A 5901");		//(= P2_P1_P3_EAX    (bv-add P2_P1_P3_EAX  0b00000000000000000000000000000001))) ;5901
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5902");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5902
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5903");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5903
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5904");		//(= P2_P1_P3_Flush    0b0)) ;5904
                                    P2_P1_P3_More = 1'b0; $display(";A 5905");		//(= P2_P1_P3_More    0b0)) ;5905
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 5906");		//(= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr )   0b01000011)) ;5906
                                    P2_P1_P3_EBX <= #1 (P2_P1_P3_EBX + 32'sb00000000000000000000000000000001); $display(";A 5907");		//(= P2_P1_P3_EBX    (bv-add P2_P1_P3_EBX  0b00000000000000000000000000000001))) ;5907
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5908");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5908
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5909");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5909
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5910");		//(= P2_P1_P3_Flush    0b0)) ;5910
                                    P2_P1_P3_More = 1'b0; $display(";A 5911");		//(= P2_P1_P3_More    0b0)) ;5911
                                end
                            default:
                                begin
                                    $display(";A 5912");		//(= (and (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b10010000) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b01100110) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b11101011) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b11101001) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b11101010) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b10110000) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b10111000) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b10111011) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b10001011) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b10001001) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b11100100) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b11100110) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b00000100) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b00000101) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b11010000) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b11000000) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b01000000) (/= ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ) 0b01000011))   true)) ;5912
                                    P2_P1_P3_InstAddrPointer = (P2_P1_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 5913");		//(= P2_P1_P3_InstAddrPointer    (bv-add P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;5913
                                    P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5914");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5914
                                    P2_P1_P3_Flush = 1'b0; $display(";A 5915");		//(= P2_P1_P3_Flush    0b0)) ;5915
                                    P2_P1_P3_More = 1'b0; $display(";A 5916");		//(= P2_P1_P3_More    0b0)) ;5916
                                end
                        endcase
                        if (((~(P2_P1_P3_InstQueueRd_Addr < P2_P1_P3_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P2_P1_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P2_P1_P3_Flush) | P2_P1_P3_More))) begin
                            $display(";A 5917");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P1_P3_InstQueueRd_Addr  P2_P1_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P1_P3_Flush ) P2_P1_P3_More ))   0b1)) ;5917
                            P2_P1_P3_State2 = 4'sb0111; $display(";A 5919");		//(= P2_P1_P3_State2    0b0111)) ;5919
                        end
                        else begin
                            $display(";A 5918");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P1_P3_InstQueueRd_Addr  P2_P1_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P1_P3_Flush ) P2_P1_P3_More ))   0b0)) ;5918
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 5920");		//(= P2_P1_P3_State2    0b0110)) ;5920
                        P2_P1_P3_Datao <= #1 ((P2_P1_P3_uWord * 32'b00000000000000010000000000000000) + P2_P1_P3_lWord); $display(";A 5921");		//(= P2_P1_P3_Datao    (bv-add (bv-mul P2_P1_P3_uWord  0b00000000000000010000000000000000) P2_P1_P3_lWord ))) ;5921
                        if ((P2_P1_P3_READY_n == 1'b0)) begin
                            $display(";A 5922");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b1)) ;5922
                            P2_P1_P3_RequestPending <= #1 1'b0; $display(";A 5924");		//(= P2_P1_P3_RequestPending    0b0)) ;5924
                            P2_P1_P3_State2 = 4'sb0101; $display(";A 5925");		//(= P2_P1_P3_State2    0b0101)) ;5925
                        end
                        else begin
                            $display(";A 5923");		//(= (bv-comp P2_P1_P3_READY_n  0b0)   0b0)) ;5923
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 5926");		//(= P2_P1_P3_State2    0b0111)) ;5926
                        if (P2_P1_P3_Flush) begin
                            $display(";A 5927");		//(= P2_P1_P3_Flush    0b1)) ;5927
                            P2_P1_P3_InstQueueRd_Addr = 5'sb00001; $display(";A 5929");		//(= P2_P1_P3_InstQueueRd_Addr    0b00001)) ;5929
                            P2_P1_P3_InstQueueWr_Addr = 5'sb00001; $display(";A 5930");		//(= P2_P1_P3_InstQueueWr_Addr    0b00001)) ;5930
                            if ((P2_P1_P3_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 5931");		//(= (bool-to-bv (bv-slt P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;5931
                                P2_P1_P3_fWord = (-P2_P1_P3_InstAddrPointer); $display(";A 5933");		//(= P2_P1_P3_fWord    (bv-neg P2_P1_P3_InstAddrPointer ))) ;5933
                            end
                            else begin
                                $display(";A 5932");		//(= (bool-to-bv (bv-slt P2_P1_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;5932
                                P2_P1_P3_fWord = P2_P1_P3_InstAddrPointer; $display(";A 5934");		//(= P2_P1_P3_fWord    P2_P1_P3_InstAddrPointer )) ;5934
                            end
                            if (((P2_P1_P3_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 5935");		//(= (bv-comp (bv-smod P2_P1_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;5935
                                P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + (P2_P1_P3_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 5937");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  (bv-smod P2_P1_P3_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;5937
                            end
                            else begin
                                $display(";A 5936");		//(= (bv-comp (bv-smod P2_P1_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;5936
                            end
                        end
                        else begin
                            $display(";A 5928");		//(= P2_P1_P3_Flush    0b0)) ;5928
                        end
                        if (((32'b00000000000000000000000000001111 - P2_P1_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 5938");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;5938
                            P2_P1_P3_State2 = 4'sb1000; $display(";A 5940");		//(= P2_P1_P3_State2    0b1000)) ;5940
                            P2_P1_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 5941");		//(= P2_P1_P3_InstQueueWr_Addr    0b00000)) ;5941
                        end
                        else begin
                            $display(";A 5939");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P1_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;5939
                            P2_P1_P3_State2 = 4'sb1001; $display(";A 5942");		//(= P2_P1_P3_State2    0b1001)) ;5942
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 5943");		//(= P2_P1_P3_State2    0b1000)) ;5943
                        if ((P2_P1_P3_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 5944");		//(= (bool-to-bv (bv-le P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;5944
                            P2_P1_P3_InstQueue[P2_P1_P3_InstQueueWr_Addr] = P2_P1_P3_InstQueue[P2_P1_P3_InstQueueRd_Addr]; $display(";A 5946");		//(= P2_P1_P3_InstQueue    ( P2_P1_P3_InstQueue P2_P1_P3_InstQueueRd_Addr ))) ;5946
                            P2_P1_P3_InstQueueRd_Addr = ((P2_P1_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5947");		//(= P2_P1_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5947
                            P2_P1_P3_InstQueueWr_Addr = ((P2_P1_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 5948");		//(= P2_P1_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P1_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;5948
                            P2_P1_P3_State2 = 4'sb1000; $display(";A 5949");		//(= P2_P1_P3_State2    0b1000)) ;5949
                        end
                        else begin
                            $display(";A 5945");		//(= (bool-to-bv (bv-le P2_P1_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;5945
                            P2_P1_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 5950");		//(= P2_P1_P3_InstQueueRd_Addr    0b00000)) ;5950
                            P2_P1_P3_State2 = 4'sb1001; $display(";A 5951");		//(= P2_P1_P3_State2    0b1001)) ;5951
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 5952");		//(= P2_P1_P3_State2    0b1001)) ;5952
                        P2_P1_P3_rEIP <= #1 P2_P1_P3_PhyAddrPointer; $display(";A 5953");		//(= P2_P1_P3_rEIP    P2_P1_P3_PhyAddrPointer )) ;5953
                        P2_P1_P3_State2 = 4'sb0001; $display(";A 5954");		//(= P2_P1_P3_State2    0b0001)) ;5954
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9016
    always @(posedge P2_P1_P3_RESET or posedge P2_P1_P3_CLOCK) begin
        if ((P2_P1_P3_RESET == 1'b1)) begin
            $display(";A 5955");		//(= (bv-comp P2_P1_P3_RESET  0b1)   0b1)) ;5955
            P2_P1_P3_ByteEnable <= #1 4'b0000; $display(";A 5957");		//(= P2_P1_P3_ByteEnable    0b0000)) ;5957
            P2_P1_P3_NonAligned <= #1 1'b0; $display(";A 5958");		//(= P2_P1_P3_NonAligned    0b0)) ;5958
        end
        else begin
            $display(";A 5956");		//(= (bv-comp P2_P1_P3_RESET  0b1)   0b0)) ;5956
            case (P2_P1_P3_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 5959");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000000)) ;5959
                        case ((P2_P1_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 5960");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;5960
                                    P2_P1_P3_ByteEnable <= #1 4'b1110; $display(";A 5961");		//(= P2_P1_P3_ByteEnable    0b1110)) ;5961
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 5962");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;5962
                                    P2_P1_P3_ByteEnable <= #1 4'b1101; $display(";A 5963");		//(= P2_P1_P3_ByteEnable    0b1101)) ;5963
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 5964");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;5964
                                    P2_P1_P3_ByteEnable <= #1 4'b1011; $display(";A 5965");		//(= P2_P1_P3_ByteEnable    0b1011)) ;5965
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 5966");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;5966
                                    P2_P1_P3_ByteEnable <= #1 4'b0111; $display(";A 5967");		//(= P2_P1_P3_ByteEnable    0b0111)) ;5967
                                end
                            default:
                                begin
                                    $display(";A 5968");		//(= (and (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;5968
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 5969");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000001)) ;5969
                        case ((P2_P1_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 5970");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;5970
                                    P2_P1_P3_ByteEnable <= #1 4'b1100; $display(";A 5971");		//(= P2_P1_P3_ByteEnable    0b1100)) ;5971
                                    P2_P1_P3_NonAligned <= #1 1'b0; $display(";A 5972");		//(= P2_P1_P3_NonAligned    0b0)) ;5972
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 5973");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;5973
                                    P2_P1_P3_ByteEnable <= #1 4'b1001; $display(";A 5974");		//(= P2_P1_P3_ByteEnable    0b1001)) ;5974
                                    P2_P1_P3_NonAligned <= #1 1'b0; $display(";A 5975");		//(= P2_P1_P3_NonAligned    0b0)) ;5975
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 5976");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;5976
                                    P2_P1_P3_ByteEnable <= #1 4'b0011; $display(";A 5977");		//(= P2_P1_P3_ByteEnable    0b0011)) ;5977
                                    P2_P1_P3_NonAligned <= #1 1'b0; $display(";A 5978");		//(= P2_P1_P3_NonAligned    0b0)) ;5978
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 5979");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;5979
                                    P2_P1_P3_ByteEnable <= #1 4'b0111; $display(";A 5980");		//(= P2_P1_P3_ByteEnable    0b0111)) ;5980
                                    P2_P1_P3_NonAligned <= #1 1'b1; $display(";A 5981");		//(= P2_P1_P3_NonAligned    0b1)) ;5981
                                end
                            default:
                                begin
                                    $display(";A 5982");		//(= (and (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;5982
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 5983");		//(= P2_P1_P3_DataWidth    0b00000000000000000000000000000010)) ;5983
                        case ((P2_P1_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 5984");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;5984
                                    P2_P1_P3_ByteEnable <= #1 4'b0000; $display(";A 5985");		//(= P2_P1_P3_ByteEnable    0b0000)) ;5985
                                    P2_P1_P3_NonAligned <= #1 1'b0; $display(";A 5986");		//(= P2_P1_P3_NonAligned    0b0)) ;5986
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 5987");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;5987
                                    P2_P1_P3_ByteEnable <= #1 4'b0001; $display(";A 5988");		//(= P2_P1_P3_ByteEnable    0b0001)) ;5988
                                    P2_P1_P3_NonAligned <= #1 1'b1; $display(";A 5989");		//(= P2_P1_P3_NonAligned    0b1)) ;5989
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 5990");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;5990
                                    P2_P1_P3_NonAligned <= #1 1'b1; $display(";A 5991");		//(= P2_P1_P3_NonAligned    0b1)) ;5991
                                    P2_P1_P3_ByteEnable <= #1 4'b0011; $display(";A 5992");		//(= P2_P1_P3_ByteEnable    0b0011)) ;5992
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 5993");		//(= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;5993
                                    P2_P1_P3_NonAligned <= #1 1'b1; $display(";A 5994");		//(= P2_P1_P3_NonAligned    0b1)) ;5994
                                    P2_P1_P3_ByteEnable <= #1 4'b0111; $display(";A 5995");		//(= P2_P1_P3_ByteEnable    0b0111)) ;5995
                                end
                            default:
                                begin
                                    $display(";A 5996");		//(= (and (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P1_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;5996
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 5997");		//(= (and (/= P2_P1_P3_DataWidth  0b00000000000000000000000000000000) (/= P2_P1_P3_DataWidth  0b00000000000000000000000000000001) (/= P2_P1_P3_DataWidth  0b00000000000000000000000000000010))   true)) ;5997
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9162
    always @(posedge P2_P2_reset or posedge P2_P2_clock) begin
        if ((P2_P2_reset == 1'b1)) begin
            P2_P2_buf1 <= #1 32'sb00000000000000000000000000000000; $display(";A 6000");		//(= P2_P2_buf1    0b00000000000000000000000000000000)) ;6000
            P2_P2_ready11 <= #1 1'b0; $display(";A 6001");		//(= P2_P2_ready11    0b0)) ;6001
            P2_P2_ready12 <= #1 1'b0; $display(";A 6002");		//(= P2_P2_ready12    0b0)) ;6002
        end
        else begin
            if (((((((P2_P2_addr1 > 30'b100000000000000000000000000000) & (P2_P2_ads1 == 1'b0)) & (P2_P2_mio1 == 1'b1)) & (P2_P2_dc1 == 1'b0)) & (P2_P2_wr1 == 1'b1)) & (P2_P2_be1 == 4'b0000))) begin
                $display(";A 6003");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P2_addr1  0b100000000000000000000000000000)) (bv-comp P2_P2_ads1  0b0)) (bv-comp P2_P2_mio1  0b1)) (bv-comp P2_P2_dc1  0b0)) (bv-comp P2_P2_wr1  0b1)) (bv-comp P2_P2_be1  0b0000))   0b1)) ;6003
                P2_P2_buf1 <= #1 P2_P2_do1; $display(";A 6005");		//(= P2_P2_buf1    P2_P2_do1 )) ;6005
                P2_P2_ready11 <= #1 1'b0; $display(";A 6006");		//(= P2_P2_ready11    0b0)) ;6006
                P2_P2_ready12 <= #1 1'b1; $display(";A 6007");		//(= P2_P2_ready12    0b1)) ;6007
            end
            else begin
                $display(";A 6004");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P2_addr1  0b100000000000000000000000000000)) (bv-comp P2_P2_ads1  0b0)) (bv-comp P2_P2_mio1  0b1)) (bv-comp P2_P2_dc1  0b0)) (bv-comp P2_P2_wr1  0b1)) (bv-comp P2_P2_be1  0b0000))   0b0)) ;6004
                if (((((((P2_P2_addr2 > 30'b100000000000000000000000000000) & (P2_P2_ads2 == 1'b0)) & (P2_P2_mio2 == 1'b1)) & (P2_P2_dc2 == 1'b0)) & (P2_P2_wr2 == 1'b1)) & (P2_P2_be2 == 4'b0000))) begin
                    $display(";A 6008");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P2_addr2  0b100000000000000000000000000000)) (bv-comp P2_P2_ads2  0b0)) (bv-comp P2_P2_mio2  0b1)) (bv-comp P2_P2_dc2  0b0)) (bv-comp P2_P2_wr2  0b1)) (bv-comp P2_P2_be2  0b0000))   0b1)) ;6008
                    P2_P2_buf1 <= #1 P2_P2_do2; $display(";A 6010");		//(= P2_P2_buf1    P2_P2_do2 )) ;6010
                    P2_P2_ready11 <= #1 1'b1; $display(";A 6011");		//(= P2_P2_ready11    0b1)) ;6011
                    P2_P2_ready12 <= #1 1'b0; $display(";A 6012");		//(= P2_P2_ready12    0b0)) ;6012
                end
                else begin
                    $display(";A 6009");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-gt P2_P2_addr2  0b100000000000000000000000000000)) (bv-comp P2_P2_ads2  0b0)) (bv-comp P2_P2_mio2  0b1)) (bv-comp P2_P2_dc2  0b0)) (bv-comp P2_P2_wr2  0b1)) (bv-comp P2_P2_be2  0b0000))   0b0)) ;6009
                    P2_P2_ready11 <= #1 1'b1; $display(";A 6013");		//(= P2_P2_ready11    0b1)) ;6013
                    P2_P2_ready12 <= #1 1'b1; $display(";A 6014");		//(= P2_P2_ready12    0b1)) ;6014
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9191
    always @(posedge P2_P2_reset or posedge P2_P2_clock) begin
        if ((P2_P2_reset == 1'b1)) begin
            P2_P2_buf2 <= #1 32'sb00000000000000000000000000000000; $display(";A 6017");		//(= P2_P2_buf2    0b00000000000000000000000000000000)) ;6017
            P2_P2_ready21 <= #1 1'b0; $display(";A 6018");		//(= P2_P2_ready21    0b0)) ;6018
            P2_P2_ready22 <= #1 1'b0; $display(";A 6019");		//(= P2_P2_ready22    0b0)) ;6019
        end
        else begin
            if (((((((P2_P2_addr2 < 30'b100000000000000000000000000000) & (P2_P2_ads2 == 1'b0)) & (P2_P2_mio2 == 1'b1)) & (P2_P2_dc2 == 1'b0)) & (P2_P2_wr2 == 1'b1)) & (P2_P2_be2 == 4'b0000))) begin
                $display(";A 6020");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P2_P2_addr2  0b100000000000000000000000000000)) (bv-comp P2_P2_ads2  0b0)) (bv-comp P2_P2_mio2  0b1)) (bv-comp P2_P2_dc2  0b0)) (bv-comp P2_P2_wr2  0b1)) (bv-comp P2_P2_be2  0b0000))   0b1)) ;6020
                P2_P2_buf2 <= #1 P2_P2_do2; $display(";A 6022");		//(= P2_P2_buf2    P2_P2_do2 )) ;6022
                P2_P2_ready21 <= #1 1'b0; $display(";A 6023");		//(= P2_P2_ready21    0b0)) ;6023
                P2_P2_ready22 <= #1 1'b1; $display(";A 6024");		//(= P2_P2_ready22    0b1)) ;6024
            end
            else begin
                $display(";A 6021");		//(= (bv-and (bv-and (bv-and (bv-and (bv-and (bool-to-bv (bv-lt P2_P2_addr2  0b100000000000000000000000000000)) (bv-comp P2_P2_ads2  0b0)) (bv-comp P2_P2_mio2  0b1)) (bv-comp P2_P2_dc2  0b0)) (bv-comp P2_P2_wr2  0b1)) (bv-comp P2_P2_be2  0b0000))   0b0)) ;6021
                if ((((((P2_P2_ads3 == 1'b0) & (P2_P2_mio3 == 1'b1)) & (P2_P2_dc3 == 1'b0)) & (P2_P2_wr3 == 1'b0)) & (P2_P2_be3 == 4'b0000))) begin
                    $display(";A 6025");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P2_P2_ads3  0b0) (bv-comp P2_P2_mio3  0b1)) (bv-comp P2_P2_dc3  0b0)) (bv-comp P2_P2_wr3  0b0)) (bv-comp P2_P2_be3  0b0000))   0b1)) ;6025
                    P2_P2_ready21 <= #1 1'b1; $display(";A 6027");		//(= P2_P2_ready21    0b1)) ;6027
                    P2_P2_ready22 <= #1 1'b0; $display(";A 6028");		//(= P2_P2_ready22    0b0)) ;6028
                end
                else begin
                    $display(";A 6026");		//(= (bv-and (bv-and (bv-and (bv-and (bv-comp P2_P2_ads3  0b0) (bv-comp P2_P2_mio3  0b1)) (bv-comp P2_P2_dc3  0b0)) (bv-comp P2_P2_wr3  0b0)) (bv-comp P2_P2_be3  0b0000))   0b0)) ;6026
                    P2_P2_ready21 <= #1 1'b1; $display(";A 6029");		//(= P2_P2_ready21    0b1)) ;6029
                    P2_P2_ready22 <= #1 1'b1; $display(";A 6030");		//(= P2_P2_ready22    0b1)) ;6030
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9219
    always @(P2_P2_datai or P2_P2_buf1 or P2_P2_addr1) begin
        if ((P2_P2_addr1 > 30'b100000000000000000000000000000)) begin
            $display(";A 6031");		//(= (bool-to-bv (bv-gt P2_P2_addr1  0b100000000000000000000000000000))   0b1)) ;6031
            P2_P2_di1 <= #1 P2_P2_buf1; $display(";A 6033");		//(= P2_P2_di1    P2_P2_buf1 )) ;6033
        end
        else begin
            $display(";A 6032");		//(= (bool-to-bv (bv-gt P2_P2_addr1  0b100000000000000000000000000000))   0b0)) ;6032
            P2_P2_di1 <= #1 P2_P2_datai; $display(";A 6034");		//(= P2_P2_di1    P2_P2_datai )) ;6034
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9225
    always @(P2_P2_buf2 or P2_P2_buf1 or P2_P2_addr2) begin
        if ((P2_P2_addr2 > 30'b100000000000000000000000000000)) begin
            $display(";A 6035");		//(= (bool-to-bv (bv-gt P2_P2_addr2  0b100000000000000000000000000000))   0b1)) ;6035
            P2_P2_di2 <= #1 P2_P2_buf1; $display(";A 6037");		//(= P2_P2_di2    P2_P2_buf1 )) ;6037
        end
        else begin
            $display(";A 6036");		//(= (bool-to-bv (bv-gt P2_P2_addr2  0b100000000000000000000000000000))   0b0)) ;6036
            P2_P2_di2 <= #1 P2_P2_buf2; $display(";A 6038");		//(= P2_P2_di2    P2_P2_buf2 )) ;6038
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9231
    always @(P2_P2_do3 or P2_P2_do2 or P2_P2_do1 or P2_P2_addr3 or P2_P2_addr2) begin
        if ((((P2_P2_do1 < 32'b00000000000000000000000000000000) & (P2_P2_do2 < 32'b00000000000000000000000000000000)) & (P2_P2_do3 < 32'b00000000000000000000000000000000))) begin
            $display(";A 6039");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P2_P2_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P2_P2_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P2_P2_do3  0b00000000000000000000000000000000)))   0b1)) ;6039
            P2_P2_address2 <= #1 P2_P2_addr3; $display(";A 6041");		//(= P2_P2_address2    P2_P2_addr3 )) ;6041
        end
        else begin
            $display(";A 6040");		//(= (bv-and (bv-and (bool-to-bv (bv-lt P2_P2_do1  0b00000000000000000000000000000000)) (bool-to-bv (bv-lt P2_P2_do2  0b00000000000000000000000000000000))) (bool-to-bv (bv-lt P2_P2_do3  0b00000000000000000000000000000000)))   0b0)) ;6040
            P2_P2_address2 <= #1 P2_P2_addr2; $display(";A 6042");		//(= P2_P2_address2    P2_P2_addr2 )) ;6042
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9237
    always @(P2_P2_ready22 or P2_P2_ready21 or P2_P2_ready12 or P2_P2_ready11 or P2_P2_ready2 or P2_P2_ready1 or P2_P2_ads3 or P2_P2_ads1 or P2_P2_mio3 or P2_P2_dc3 or P2_P2_wr3 or P2_P2_addr1 or P2_P2_do3 or P2_P2_buf2) begin
        P2_P2_di3 <= #1 P2_P2_buf2; $display(";A 6043");		//(= P2_P2_di3    P2_P2_buf2 )) ;6043
        P2_P2_datao <= #1 P2_P2_do3; $display(";A 6044");		//(= P2_P2_datao    P2_P2_do3 )) ;6044
        P2_P2_address1 <= #1 P2_P2_addr1; $display(";A 6045");		//(= P2_P2_address1    P2_P2_addr1 )) ;6045
        P2_P2_wr <= #1 P2_P2_wr3; $display(";A 6046");		//(= P2_P2_wr    P2_P2_wr3 )) ;6046
        P2_P2_dc <= #1 P2_P2_dc3; $display(";A 6047");		//(= P2_P2_dc    P2_P2_dc3 )) ;6047
        P2_P2_mio <= #1 P2_P2_mio3; $display(";A 6048");		//(= P2_P2_mio    P2_P2_mio3 )) ;6048
        P2_P2_ast1 <= #1 P2_P2_ads1; $display(";A 6049");		//(= P2_P2_ast1    P2_P2_ads1 )) ;6049
        P2_P2_ast2 <= #1 P2_P2_ads3; $display(";A 6050");		//(= P2_P2_ast2    P2_P2_ads3 )) ;6050
        P2_P2_rdy1 <= #1 (P2_P2_ready11 & P2_P2_ready1); $display(";A 6051");		//(= P2_P2_rdy1    (bv-and P2_P2_ready11  P2_P2_ready1 ))) ;6051
        P2_P2_rdy2 <= #1 (P2_P2_ready12 & P2_P2_ready21); $display(";A 6052");		//(= P2_P2_rdy2    (bv-and P2_P2_ready12  P2_P2_ready21 ))) ;6052
        P2_P2_rdy3 <= #1 (P2_P2_ready22 & P2_P2_ready2); $display(";A 6053");		//(= P2_P2_rdy3    (bv-and P2_P2_ready22  P2_P2_ready2 ))) ;6053
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9362
    always @(posedge P2_P2_P1_RESET or posedge P2_P2_P1_CLOCK) begin
        if ((P2_P2_P1_RESET == 1'b1)) begin
            $display(";A 6054");		//(= (bv-comp P2_P2_P1_RESET  0b1)   0b1)) ;6054
            P2_P2_P1_BE_n <= #1 4'b0000; $display(";A 6056");		//(= P2_P2_P1_BE_n    0b0000)) ;6056
            P2_P2_P1_Address <= #1 30'sb000000000000000000000000000000; $display(";A 6057");		//(= P2_P2_P1_Address    0b000000000000000000000000000000)) ;6057
            P2_P2_P1_W_R_n <= #1 1'b0; $display(";A 6058");		//(= P2_P2_P1_W_R_n    0b0)) ;6058
            P2_P2_P1_D_C_n <= #1 1'b0; $display(";A 6059");		//(= P2_P2_P1_D_C_n    0b0)) ;6059
            P2_P2_P1_M_IO_n <= #1 1'b0; $display(";A 6060");		//(= P2_P2_P1_M_IO_n    0b0)) ;6060
            P2_P2_P1_ADS_n <= #1 1'b0; $display(";A 6061");		//(= P2_P2_P1_ADS_n    0b0)) ;6061
            P2_P2_P1_State <= #1 3'sb000; $display(";A 6062");		//(= P2_P2_P1_State    0b000)) ;6062
            P2_P2_P1_StateNA <= #1 1'b0; $display(";A 6063");		//(= P2_P2_P1_StateNA    0b0)) ;6063
            P2_P2_P1_StateBS16 <= #1 1'b0; $display(";A 6064");		//(= P2_P2_P1_StateBS16    0b0)) ;6064
            P2_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 6065");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000000)) ;6065
        end
        else begin
            $display(";A 6055");		//(= (bv-comp P2_P2_P1_RESET  0b1)   0b0)) ;6055
            case (P2_P2_P1_State)
                3'b000 :
                    begin
                        $display(";A 6066");		//(= P2_P2_P1_State    0b000)) ;6066
                        P2_P2_P1_D_C_n <= #1 1'b1; $display(";A 6067");		//(= P2_P2_P1_D_C_n    0b1)) ;6067
                        P2_P2_P1_ADS_n <= #1 1'b1; $display(";A 6068");		//(= P2_P2_P1_ADS_n    0b1)) ;6068
                        P2_P2_P1_State <= #1 3'sb001; $display(";A 6069");		//(= P2_P2_P1_State    0b001)) ;6069
                        P2_P2_P1_StateNA <= #1 1'b1; $display(";A 6070");		//(= P2_P2_P1_StateNA    0b1)) ;6070
                        P2_P2_P1_StateBS16 <= #1 1'b1; $display(";A 6071");		//(= P2_P2_P1_StateBS16    0b1)) ;6071
                        P2_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 6072");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;6072
                        P2_P2_P1_State <= #1 3'sb001; $display(";A 6073");		//(= P2_P2_P1_State    0b001)) ;6073
                    end
                3'b001 :
                    begin
                        $display(";A 6074");		//(= P2_P2_P1_State    0b001)) ;6074
                        if ((P2_P2_P1_RequestPending == 1'b1)) begin
                            $display(";A 6075");		//(= (bv-comp P2_P2_P1_RequestPending  0b1)   0b1)) ;6075
                            P2_P2_P1_State <= #1 3'sb010; $display(";A 6077");		//(= P2_P2_P1_State    0b010)) ;6077
                        end
                        else begin
                            $display(";A 6076");		//(= (bv-comp P2_P2_P1_RequestPending  0b1)   0b0)) ;6076
                            if ((P2_P2_P1_HOLD == 1'b1)) begin
                                $display(";A 6078");		//(= (bv-comp P2_P2_P1_HOLD  0b1)   0b1)) ;6078
                                P2_P2_P1_State <= #1 3'sb101; $display(";A 6080");		//(= P2_P2_P1_State    0b101)) ;6080
                            end
                            else begin
                                $display(";A 6079");		//(= (bv-comp P2_P2_P1_HOLD  0b1)   0b0)) ;6079
                                P2_P2_P1_State <= #1 3'sb001; $display(";A 6081");		//(= P2_P2_P1_State    0b001)) ;6081
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 6082");		//(= P2_P2_P1_State    0b010)) ;6082
                        P2_P2_P1_Address <= #1 ((P2_P2_P1_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 6083");		//(= P2_P2_P1_Address    (bv-smod (bv-sdiv P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;6083
                        P2_P2_P1_BE_n <= #1 P2_P2_P1_ByteEnable; $display(";A 6084");		//(= P2_P2_P1_BE_n    P2_P2_P1_ByteEnable )) ;6084
                        P2_P2_P1_M_IO_n <= #1 P2_P2_P1_MemoryFetch; $display(";A 6085");		//(= P2_P2_P1_M_IO_n    P2_P2_P1_MemoryFetch )) ;6085
                        if ((P2_P2_P1_ReadRequest == 1'b1)) begin
                            $display(";A 6086");		//(= (bv-comp P2_P2_P1_ReadRequest  0b1)   0b1)) ;6086
                            P2_P2_P1_W_R_n <= #1 1'b0; $display(";A 6088");		//(= P2_P2_P1_W_R_n    0b0)) ;6088
                        end
                        else begin
                            $display(";A 6087");		//(= (bv-comp P2_P2_P1_ReadRequest  0b1)   0b0)) ;6087
                            P2_P2_P1_W_R_n <= #1 1'b1; $display(";A 6089");		//(= P2_P2_P1_W_R_n    0b1)) ;6089
                        end
                        if ((P2_P2_P1_CodeFetch == 1'b1)) begin
                            $display(";A 6090");		//(= (bv-comp P2_P2_P1_CodeFetch  0b1)   0b1)) ;6090
                            P2_P2_P1_D_C_n <= #1 1'b0; $display(";A 6092");		//(= P2_P2_P1_D_C_n    0b0)) ;6092
                        end
                        else begin
                            $display(";A 6091");		//(= (bv-comp P2_P2_P1_CodeFetch  0b1)   0b0)) ;6091
                            P2_P2_P1_D_C_n <= #1 1'b1; $display(";A 6093");		//(= P2_P2_P1_D_C_n    0b1)) ;6093
                        end
                        P2_P2_P1_ADS_n <= #1 1'b0; $display(";A 6094");		//(= P2_P2_P1_ADS_n    0b0)) ;6094
                        P2_P2_P1_State <= #1 3'sb011; $display(";A 6095");		//(= P2_P2_P1_State    0b011)) ;6095
                    end
                3'b011 :
                    begin
                        $display(";A 6096");		//(= P2_P2_P1_State    0b011)) ;6096
                        if ((((P2_P2_P1_READY_n == 1'b0) & (P2_P2_P1_HOLD == 1'b0)) & (P2_P2_P1_RequestPending == 1'b1))) begin
                            $display(";A 6097");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b1))   0b1)) ;6097
                            P2_P2_P1_State <= #1 3'sb010; $display(";A 6099");		//(= P2_P2_P1_State    0b010)) ;6099
                        end
                        else begin
                            $display(";A 6098");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b1))   0b0)) ;6098
                            if (((P2_P2_P1_READY_n == 1'b1) & (P2_P2_P1_NA_n == 1'b1))) begin
                                $display(";A 6100");		//(= (bv-and (bv-comp P2_P2_P1_READY_n  0b1) (bv-comp P2_P2_P1_NA_n  0b1))   0b1)) ;6100
                            end
                            else begin
                                $display(";A 6101");		//(= (bv-and (bv-comp P2_P2_P1_READY_n  0b1) (bv-comp P2_P2_P1_NA_n  0b1))   0b0)) ;6101
                                if ((((P2_P2_P1_RequestPending == 1'b1) | (P2_P2_P1_HOLD == 1'b1)) & ((P2_P2_P1_READY_n == 1'b1) & (P2_P2_P1_NA_n == 1'b0)))) begin
                                    $display(";A 6102");		//(= (bv-and (bv-or (bv-comp P2_P2_P1_RequestPending  0b1) (bv-comp P2_P2_P1_HOLD  0b1)) (bv-and (bv-comp P2_P2_P1_READY_n  0b1) (bv-comp P2_P2_P1_NA_n  0b0)))   0b1)) ;6102
                                    P2_P2_P1_State <= #1 3'sb111; $display(";A 6104");		//(= P2_P2_P1_State    0b111)) ;6104
                                end
                                else begin
                                    $display(";A 6103");		//(= (bv-and (bv-or (bv-comp P2_P2_P1_RequestPending  0b1) (bv-comp P2_P2_P1_HOLD  0b1)) (bv-and (bv-comp P2_P2_P1_READY_n  0b1) (bv-comp P2_P2_P1_NA_n  0b0)))   0b0)) ;6103
                                    if (((((P2_P2_P1_RequestPending == 1'b1) & (P2_P2_P1_HOLD == 1'b0)) & (P2_P2_P1_READY_n == 1'b1)) & (P2_P2_P1_NA_n == 1'b0))) begin
                                        $display(";A 6105");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P2_P1_RequestPending  0b1) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_READY_n  0b1)) (bv-comp P2_P2_P1_NA_n  0b0))   0b1)) ;6105
                                        P2_P2_P1_State <= #1 3'sb110; $display(";A 6107");		//(= P2_P2_P1_State    0b110)) ;6107
                                    end
                                    else begin
                                        $display(";A 6106");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P2_P1_RequestPending  0b1) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_READY_n  0b1)) (bv-comp P2_P2_P1_NA_n  0b0))   0b0)) ;6106
                                        if ((((P2_P2_P1_RequestPending == 1'b0) & (P2_P2_P1_HOLD == 1'b0)) & (P2_P2_P1_READY_n == 1'b0))) begin
                                            $display(";A 6108");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_RequestPending  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_READY_n  0b0))   0b1)) ;6108
                                            P2_P2_P1_State <= #1 3'sb001; $display(";A 6110");		//(= P2_P2_P1_State    0b001)) ;6110
                                        end
                                        else begin
                                            $display(";A 6109");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_RequestPending  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_READY_n  0b0))   0b0)) ;6109
                                            if (((P2_P2_P1_HOLD == 1'b1) & (P2_P2_P1_READY_n == 1'b1))) begin
                                                $display(";A 6111");		//(= (bv-and (bv-comp P2_P2_P1_HOLD  0b1) (bv-comp P2_P2_P1_READY_n  0b1))   0b1)) ;6111
                                                P2_P2_P1_State <= #1 3'sb101; $display(";A 6113");		//(= P2_P2_P1_State    0b101)) ;6113
                                            end
                                            else begin
                                                $display(";A 6112");		//(= (bv-and (bv-comp P2_P2_P1_HOLD  0b1) (bv-comp P2_P2_P1_READY_n  0b1))   0b0)) ;6112
                                                P2_P2_P1_State <= #1 3'sb011; $display(";A 6114");		//(= P2_P2_P1_State    0b011)) ;6114
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P2_P2_P1_StateBS16 <= #1 P2_P2_P1_BS16_n; $display(";A 6115");		//(= P2_P2_P1_StateBS16    P2_P2_P1_BS16_n )) ;6115
                        if ((P2_P2_P1_BS16_n == 1'b0)) begin
                            $display(";A 6116");		//(= (bv-comp P2_P2_P1_BS16_n  0b0)   0b1)) ;6116
                            P2_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 6118");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000001)) ;6118
                        end
                        else begin
                            $display(";A 6117");		//(= (bv-comp P2_P2_P1_BS16_n  0b0)   0b0)) ;6117
                            P2_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 6119");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;6119
                        end
                        P2_P2_P1_StateNA <= #1 P2_P2_P1_NA_n; $display(";A 6120");		//(= P2_P2_P1_StateNA    P2_P2_P1_NA_n )) ;6120
                        P2_P2_P1_ADS_n <= #1 1'b1; $display(";A 6121");		//(= P2_P2_P1_ADS_n    0b1)) ;6121
                    end
                3'b100 :
                    begin
                        $display(";A 6122");		//(= P2_P2_P1_State    0b100)) ;6122
                        if ((((P2_P2_P1_NA_n == 1'b0) & (P2_P2_P1_HOLD == 1'b0)) & (P2_P2_P1_RequestPending == 1'b1))) begin
                            $display(";A 6123");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_NA_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b1))   0b1)) ;6123
                            P2_P2_P1_State <= #1 3'sb110; $display(";A 6125");		//(= P2_P2_P1_State    0b110)) ;6125
                        end
                        else begin
                            $display(";A 6124");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_NA_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b1))   0b0)) ;6124
                            if (((P2_P2_P1_NA_n == 1'b0) & ((P2_P2_P1_HOLD == 1'b1) | (P2_P2_P1_RequestPending == 1'b0)))) begin
                                $display(";A 6126");		//(= (bv-and (bv-comp P2_P2_P1_NA_n  0b0) (bv-or (bv-comp P2_P2_P1_HOLD  0b1) (bv-comp P2_P2_P1_RequestPending  0b0)))   0b1)) ;6126
                                P2_P2_P1_State <= #1 3'sb111; $display(";A 6128");		//(= P2_P2_P1_State    0b111)) ;6128
                            end
                            else begin
                                $display(";A 6127");		//(= (bv-and (bv-comp P2_P2_P1_NA_n  0b0) (bv-or (bv-comp P2_P2_P1_HOLD  0b1) (bv-comp P2_P2_P1_RequestPending  0b0)))   0b0)) ;6127
                                if ((P2_P2_P1_NA_n == 1'b1)) begin
                                    $display(";A 6129");		//(= (bv-comp P2_P2_P1_NA_n  0b1)   0b1)) ;6129
                                    P2_P2_P1_State <= #1 3'sb011; $display(";A 6131");		//(= P2_P2_P1_State    0b011)) ;6131
                                end
                                else begin
                                    $display(";A 6130");		//(= (bv-comp P2_P2_P1_NA_n  0b1)   0b0)) ;6130
                                    P2_P2_P1_State <= #1 3'sb100; $display(";A 6132");		//(= P2_P2_P1_State    0b100)) ;6132
                                end
                            end
                        end
                        P2_P2_P1_StateBS16 <= #1 P2_P2_P1_BS16_n; $display(";A 6133");		//(= P2_P2_P1_StateBS16    P2_P2_P1_BS16_n )) ;6133
                        if ((P2_P2_P1_BS16_n == 1'b0)) begin
                            $display(";A 6134");		//(= (bv-comp P2_P2_P1_BS16_n  0b0)   0b1)) ;6134
                            P2_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 6136");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000001)) ;6136
                        end
                        else begin
                            $display(";A 6135");		//(= (bv-comp P2_P2_P1_BS16_n  0b0)   0b0)) ;6135
                            P2_P2_P1_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 6137");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;6137
                        end
                        P2_P2_P1_StateNA <= #1 P2_P2_P1_NA_n; $display(";A 6138");		//(= P2_P2_P1_StateNA    P2_P2_P1_NA_n )) ;6138
                        P2_P2_P1_ADS_n <= #1 1'b1; $display(";A 6139");		//(= P2_P2_P1_ADS_n    0b1)) ;6139
                    end
                3'b101 :
                    begin
                        $display(";A 6140");		//(= P2_P2_P1_State    0b101)) ;6140
                        if (((P2_P2_P1_HOLD == 1'b0) & (P2_P2_P1_RequestPending == 1'b1))) begin
                            $display(";A 6141");		//(= (bv-and (bv-comp P2_P2_P1_HOLD  0b0) (bv-comp P2_P2_P1_RequestPending  0b1))   0b1)) ;6141
                            P2_P2_P1_State <= #1 3'sb010; $display(";A 6143");		//(= P2_P2_P1_State    0b010)) ;6143
                        end
                        else begin
                            $display(";A 6142");		//(= (bv-and (bv-comp P2_P2_P1_HOLD  0b0) (bv-comp P2_P2_P1_RequestPending  0b1))   0b0)) ;6142
                            if (((P2_P2_P1_HOLD == 1'b0) & (P2_P2_P1_RequestPending == 1'b0))) begin
                                $display(";A 6144");		//(= (bv-and (bv-comp P2_P2_P1_HOLD  0b0) (bv-comp P2_P2_P1_RequestPending  0b0))   0b1)) ;6144
                                P2_P2_P1_State <= #1 3'sb001; $display(";A 6146");		//(= P2_P2_P1_State    0b001)) ;6146
                            end
                            else begin
                                $display(";A 6145");		//(= (bv-and (bv-comp P2_P2_P1_HOLD  0b0) (bv-comp P2_P2_P1_RequestPending  0b0))   0b0)) ;6145
                                P2_P2_P1_State <= #1 3'sb101; $display(";A 6147");		//(= P2_P2_P1_State    0b101)) ;6147
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 6148");		//(= P2_P2_P1_State    0b110)) ;6148
                        P2_P2_P1_Address <= #1 ((P2_P2_P1_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 6149");		//(= P2_P2_P1_Address    (bv-smod (bv-sdiv P2_P2_P1_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;6149
                        P2_P2_P1_BE_n <= #1 P2_P2_P1_ByteEnable; $display(";A 6150");		//(= P2_P2_P1_BE_n    P2_P2_P1_ByteEnable )) ;6150
                        P2_P2_P1_M_IO_n <= #1 P2_P2_P1_MemoryFetch; $display(";A 6151");		//(= P2_P2_P1_M_IO_n    P2_P2_P1_MemoryFetch )) ;6151
                        if ((P2_P2_P1_ReadRequest == 1'b1)) begin
                            $display(";A 6152");		//(= (bv-comp P2_P2_P1_ReadRequest  0b1)   0b1)) ;6152
                            P2_P2_P1_W_R_n <= #1 1'b0; $display(";A 6154");		//(= P2_P2_P1_W_R_n    0b0)) ;6154
                        end
                        else begin
                            $display(";A 6153");		//(= (bv-comp P2_P2_P1_ReadRequest  0b1)   0b0)) ;6153
                            P2_P2_P1_W_R_n <= #1 1'b1; $display(";A 6155");		//(= P2_P2_P1_W_R_n    0b1)) ;6155
                        end
                        if ((P2_P2_P1_CodeFetch == 1'b1)) begin
                            $display(";A 6156");		//(= (bv-comp P2_P2_P1_CodeFetch  0b1)   0b1)) ;6156
                            P2_P2_P1_D_C_n <= #1 1'b0; $display(";A 6158");		//(= P2_P2_P1_D_C_n    0b0)) ;6158
                        end
                        else begin
                            $display(";A 6157");		//(= (bv-comp P2_P2_P1_CodeFetch  0b1)   0b0)) ;6157
                            P2_P2_P1_D_C_n <= #1 1'b1; $display(";A 6159");		//(= P2_P2_P1_D_C_n    0b1)) ;6159
                        end
                        P2_P2_P1_ADS_n <= #1 1'b0; $display(";A 6160");		//(= P2_P2_P1_ADS_n    0b0)) ;6160
                        if ((P2_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 6161");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6161
                            P2_P2_P1_State <= #1 3'sb100; $display(";A 6163");		//(= P2_P2_P1_State    0b100)) ;6163
                        end
                        else begin
                            $display(";A 6162");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6162
                            P2_P2_P1_State <= #1 3'sb110; $display(";A 6164");		//(= P2_P2_P1_State    0b110)) ;6164
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 6165");		//(= P2_P2_P1_State    0b111)) ;6165
                        if ((((P2_P2_P1_READY_n == 1'b1) & (P2_P2_P1_RequestPending == 1'b1)) & (P2_P2_P1_HOLD == 1'b0))) begin
                            $display(";A 6166");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b1) (bv-comp P2_P2_P1_RequestPending  0b1)) (bv-comp P2_P2_P1_HOLD  0b0))   0b1)) ;6166
                            P2_P2_P1_State <= #1 3'sb110; $display(";A 6168");		//(= P2_P2_P1_State    0b110)) ;6168
                        end
                        else begin
                            $display(";A 6167");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b1) (bv-comp P2_P2_P1_RequestPending  0b1)) (bv-comp P2_P2_P1_HOLD  0b0))   0b0)) ;6167
                            if (((P2_P2_P1_READY_n == 1'b0) & (P2_P2_P1_HOLD == 1'b1))) begin
                                $display(";A 6169");		//(= (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b1))   0b1)) ;6169
                                P2_P2_P1_State <= #1 3'sb101; $display(";A 6171");		//(= P2_P2_P1_State    0b101)) ;6171
                            end
                            else begin
                                $display(";A 6170");		//(= (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b1))   0b0)) ;6170
                                if ((((P2_P2_P1_READY_n == 1'b0) & (P2_P2_P1_HOLD == 1'b0)) & (P2_P2_P1_RequestPending == 1'b1))) begin
                                    $display(";A 6172");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b1))   0b1)) ;6172
                                    P2_P2_P1_State <= #1 3'sb010; $display(";A 6174");		//(= P2_P2_P1_State    0b010)) ;6174
                                end
                                else begin
                                    $display(";A 6173");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b1))   0b0)) ;6173
                                    if ((((P2_P2_P1_READY_n == 1'b0) & (P2_P2_P1_HOLD == 1'b0)) & (P2_P2_P1_RequestPending == 1'b0))) begin
                                        $display(";A 6175");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b0))   0b1)) ;6175
                                        P2_P2_P1_State <= #1 3'sb001; $display(";A 6177");		//(= P2_P2_P1_State    0b001)) ;6177
                                    end
                                    else begin
                                        $display(";A 6176");		//(= (bv-and (bv-and (bv-comp P2_P2_P1_READY_n  0b0) (bv-comp P2_P2_P1_HOLD  0b0)) (bv-comp P2_P2_P1_RequestPending  0b0))   0b0)) ;6176
                                        P2_P2_P1_State <= #1 3'sb111; $display(";A 6178");		//(= P2_P2_P1_State    0b111)) ;6178
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9506
    always @(posedge P2_P2_P1_RESET or posedge P2_P2_P1_CLOCK) begin
        if ((P2_P2_P1_RESET == 1'b1)) begin
            $display(";A 6179");		//(= (bv-comp P2_P2_P1_RESET  0b1)   0b1)) ;6179
            P2_P2_P1_State2 = 4'sb0000; $display(";A 6181");		//(= P2_P2_P1_State2    0b0000)) ;6181
            P2_P2_P1_InstQueue[0] = 8'b00000000; $display(";A 6182");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6182
            P2_P2_P1_InstQueue[1] = 8'b00000000; $display(";A 6183");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6183
            P2_P2_P1_InstQueue[2] = 8'b00000000; $display(";A 6184");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6184
            P2_P2_P1_InstQueue[3] = 8'b00000000; $display(";A 6185");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6185
            P2_P2_P1_InstQueue[4] = 8'b00000000; $display(";A 6186");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6186
            P2_P2_P1_InstQueue[5] = 8'b00000000; $display(";A 6187");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6187
            P2_P2_P1_InstQueue[6] = 8'b00000000; $display(";A 6188");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6188
            P2_P2_P1_InstQueue[7] = 8'b00000000; $display(";A 6189");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6189
            P2_P2_P1_InstQueue[8] = 8'b00000000; $display(";A 6190");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6190
            P2_P2_P1_InstQueue[9] = 8'b00000000; $display(";A 6191");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6191
            P2_P2_P1_InstQueue[10] = 8'b00000000; $display(";A 6192");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6192
            P2_P2_P1_InstQueue[11] = 8'b00000000; $display(";A 6193");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6193
            P2_P2_P1_InstQueue[12] = 8'b00000000; $display(";A 6194");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6194
            P2_P2_P1_InstQueue[13] = 8'b00000000; $display(";A 6195");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6195
            P2_P2_P1_InstQueue[14] = 8'b00000000; $display(";A 6196");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6196
            P2_P2_P1_InstQueue[15] = 8'b00000000; $display(";A 6197");		//(= P2_P2_P1_InstQueue    0b00000000)) ;6197
            P2_P2_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 6198");		//(= P2_P2_P1_InstQueueRd_Addr    0b00000)) ;6198
            P2_P2_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 6199");		//(= P2_P2_P1_InstQueueWr_Addr    0b00000)) ;6199
            P2_P2_P1_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 6200");		//(= P2_P2_P1_InstAddrPointer    0b00000000000000000000000000000000)) ;6200
            P2_P2_P1_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 6201");		//(= P2_P2_P1_PhyAddrPointer    0b00000000000000000000000000000000)) ;6201
            P2_P2_P1_Extended = 1'b0; $display(";A 6202");		//(= P2_P2_P1_Extended    0b0)) ;6202
            P2_P2_P1_More = 1'b0; $display(";A 6203");		//(= P2_P2_P1_More    0b0)) ;6203
            P2_P2_P1_Flush = 1'b0; $display(";A 6204");		//(= P2_P2_P1_Flush    0b0)) ;6204
            P2_P2_P1_lWord = 16'sb0000000000000000; $display(";A 6205");		//(= P2_P2_P1_lWord    0b0000000000000000)) ;6205
            P2_P2_P1_uWord = 15'sb000000000000000; $display(";A 6206");		//(= P2_P2_P1_uWord    0b000000000000000)) ;6206
            P2_P2_P1_fWord = 32'sb00000000000000000000000000000000; $display(";A 6207");		//(= P2_P2_P1_fWord    0b00000000000000000000000000000000)) ;6207
            P2_P2_P1_CodeFetch <= #1 1'b0; $display(";A 6208");		//(= P2_P2_P1_CodeFetch    0b0)) ;6208
            P2_P2_P1_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 6209");		//(= P2_P2_P1_Datao    0b00000000000000000000000000000000)) ;6209
            P2_P2_P1_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 6210");		//(= P2_P2_P1_EAX    0b00000000000000000000000000000000)) ;6210
            P2_P2_P1_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 6211");		//(= P2_P2_P1_EBX    0b00000000000000000000000000000000)) ;6211
            P2_P2_P1_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 6212");		//(= P2_P2_P1_rEIP    0b00000000000000000000000000000000)) ;6212
            P2_P2_P1_ReadRequest <= #1 1'b0; $display(";A 6213");		//(= P2_P2_P1_ReadRequest    0b0)) ;6213
            P2_P2_P1_MemoryFetch <= #1 1'b0; $display(";A 6214");		//(= P2_P2_P1_MemoryFetch    0b0)) ;6214
            P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6215");		//(= P2_P2_P1_RequestPending    0b0)) ;6215
        end
        else begin
            $display(";A 6180");		//(= (bv-comp P2_P2_P1_RESET  0b1)   0b0)) ;6180
            case (P2_P2_P1_State2)
                4'b0000 :
                    begin
                        $display(";A 6216");		//(= P2_P2_P1_State2    0b0000)) ;6216
                        P2_P2_P1_PhyAddrPointer = P2_P2_P1_rEIP; $display(";A 6217");		//(= P2_P2_P1_PhyAddrPointer    P2_P2_P1_rEIP )) ;6217
                        P2_P2_P1_InstAddrPointer = P2_P2_P1_PhyAddrPointer; $display(";A 6218");		//(= P2_P2_P1_InstAddrPointer    P2_P2_P1_PhyAddrPointer )) ;6218
                        P2_P2_P1_State2 = 4'sb0001; $display(";A 6219");		//(= P2_P2_P1_State2    0b0001)) ;6219
                        P2_P2_P1_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 6220");		//(= P2_P2_P1_rEIP    0b00000000000011111111111111110000)) ;6220
                        P2_P2_P1_ReadRequest <= #1 1'b1; $display(";A 6221");		//(= P2_P2_P1_ReadRequest    0b1)) ;6221
                        P2_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 6222");		//(= P2_P2_P1_MemoryFetch    0b1)) ;6222
                        P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6223");		//(= P2_P2_P1_RequestPending    0b1)) ;6223
                    end
                4'b0001 :
                    begin
                        $display(";A 6224");		//(= P2_P2_P1_State2    0b0001)) ;6224
                        P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6225");		//(= P2_P2_P1_RequestPending    0b1)) ;6225
                        P2_P2_P1_ReadRequest <= #1 1'b1; $display(";A 6226");		//(= P2_P2_P1_ReadRequest    0b1)) ;6226
                        P2_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 6227");		//(= P2_P2_P1_MemoryFetch    0b1)) ;6227
                        P2_P2_P1_CodeFetch <= #1 1'b1; $display(";A 6228");		//(= P2_P2_P1_CodeFetch    0b1)) ;6228
                        if ((P2_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 6229");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6229
                            P2_P2_P1_State2 = 4'sb0010; $display(";A 6231");		//(= P2_P2_P1_State2    0b0010)) ;6231
                        end
                        else begin
                            $display(";A 6230");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6230
                            P2_P2_P1_State2 = 4'sb0001; $display(";A 6232");		//(= P2_P2_P1_State2    0b0001)) ;6232
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 6233");		//(= P2_P2_P1_State2    0b0010)) ;6233
                        P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6234");		//(= P2_P2_P1_RequestPending    0b0)) ;6234
                        P2_P2_P1_InstQueue[P2_P2_P1_InstQueueWr_Addr] = (P2_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 6235");		//(= P2_P2_P1_InstQueue    (bv-smod P2_P2_P1_Datai  0b00000000000000000000000100000000))) ;6235
                        P2_P2_P1_InstQueueWr_Addr = ((P2_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6236");		//(= P2_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6236
                        P2_P2_P1_InstQueue[P2_P2_P1_InstQueueWr_Addr] = (P2_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 6237");		//(= P2_P2_P1_InstQueue    (bv-smod P2_P2_P1_Datai  0b00000000000000000000000100000000))) ;6237
                        P2_P2_P1_InstQueueWr_Addr = ((P2_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6238");		//(= P2_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6238
                        if ((P2_P2_P1_StateBS16 == 1'b1)) begin
                            $display(";A 6239");		//(= (bv-comp P2_P2_P1_StateBS16  0b1)   0b1)) ;6239
                            P2_P2_P1_InstQueue[P2_P2_P1_InstQueueWr_Addr] = ((P2_P2_P1_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 6241");		//(= P2_P2_P1_InstQueue    (bv-smod (bv-sdiv P2_P2_P1_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;6241
                            P2_P2_P1_InstQueueWr_Addr = ((P2_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6242");		//(= P2_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6242
                            P2_P2_P1_InstQueue[P2_P2_P1_InstQueueWr_Addr] = ((P2_P2_P1_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 6243");		//(= P2_P2_P1_InstQueue    (bv-smod (bv-sdiv P2_P2_P1_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;6243
                            P2_P2_P1_InstQueueWr_Addr = ((P2_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6244");		//(= P2_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6244
                            P2_P2_P1_PhyAddrPointer = (P2_P2_P1_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 6245");		//(= P2_P2_P1_PhyAddrPointer    (bv-add P2_P2_P1_PhyAddrPointer  0b00000000000000000000000000000100))) ;6245
                            P2_P2_P1_State2 = 4'sb0101; $display(";A 6246");		//(= P2_P2_P1_State2    0b0101)) ;6246
                        end
                        else begin
                            $display(";A 6240");		//(= (bv-comp P2_P2_P1_StateBS16  0b1)   0b0)) ;6240
                            P2_P2_P1_PhyAddrPointer = (P2_P2_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6247");		//(= P2_P2_P1_PhyAddrPointer    (bv-add P2_P2_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;6247
                            if ((P2_P2_P1_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 6248");		//(= (bool-to-bv (bv-slt P2_P2_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;6248
                                P2_P2_P1_rEIP <= #1 (-P2_P2_P1_PhyAddrPointer); $display(";A 6250");		//(= P2_P2_P1_rEIP    (bv-neg P2_P2_P1_PhyAddrPointer ))) ;6250
                            end
                            else begin
                                $display(";A 6249");		//(= (bool-to-bv (bv-slt P2_P2_P1_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;6249
                                P2_P2_P1_rEIP <= #1 P2_P2_P1_PhyAddrPointer; $display(";A 6251");		//(= P2_P2_P1_rEIP    P2_P2_P1_PhyAddrPointer )) ;6251
                            end
                            P2_P2_P1_State2 = 4'sb0011; $display(";A 6252");		//(= P2_P2_P1_State2    0b0011)) ;6252
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 6253");		//(= P2_P2_P1_State2    0b0011)) ;6253
                        P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6254");		//(= P2_P2_P1_RequestPending    0b1)) ;6254
                        if ((P2_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 6255");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6255
                            P2_P2_P1_State2 = 4'sb0100; $display(";A 6257");		//(= P2_P2_P1_State2    0b0100)) ;6257
                        end
                        else begin
                            $display(";A 6256");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6256
                            P2_P2_P1_State2 = 4'sb0011; $display(";A 6258");		//(= P2_P2_P1_State2    0b0011)) ;6258
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 6259");		//(= P2_P2_P1_State2    0b0100)) ;6259
                        P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6260");		//(= P2_P2_P1_RequestPending    0b0)) ;6260
                        P2_P2_P1_InstQueue[P2_P2_P1_InstQueueWr_Addr] = (P2_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 6261");		//(= P2_P2_P1_InstQueue    (bv-smod P2_P2_P1_Datai  0b00000000000000000000000100000000))) ;6261
                        P2_P2_P1_InstQueueWr_Addr = ((P2_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6262");		//(= P2_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6262
                        P2_P2_P1_InstQueue[P2_P2_P1_InstQueueWr_Addr] = (P2_P2_P1_Datai % 32'b00000000000000000000000100000000); $display(";A 6263");		//(= P2_P2_P1_InstQueue    (bv-smod P2_P2_P1_Datai  0b00000000000000000000000100000000))) ;6263
                        P2_P2_P1_InstQueueWr_Addr = ((P2_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6264");		//(= P2_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6264
                        P2_P2_P1_PhyAddrPointer = (P2_P2_P1_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6265");		//(= P2_P2_P1_PhyAddrPointer    (bv-add P2_P2_P1_PhyAddrPointer  0b00000000000000000000000000000010))) ;6265
                        P2_P2_P1_State2 = 4'sb0101; $display(";A 6266");		//(= P2_P2_P1_State2    0b0101)) ;6266
                    end
                4'b0101 :
                    begin
                        $display(";A 6267");		//(= P2_P2_P1_State2    0b0101)) ;6267
                        case (P2_P2_P1_InstQueue[P2_P2_P1_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 6268");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b10010000)) ;6268
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6269");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6269
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6270");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6270
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6271");		//(= P2_P2_P1_Flush    0b0)) ;6271
                                    P2_P2_P1_More = 1'b0; $display(";A 6272");		//(= P2_P2_P1_More    0b0)) ;6272
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 6273");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b01100110)) ;6273
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6274");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6274
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6275");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6275
                                    P2_P2_P1_Extended = 1'b1; $display(";A 6276");		//(= P2_P2_P1_Extended    0b1)) ;6276
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6277");		//(= P2_P2_P1_Flush    0b0)) ;6277
                                    P2_P2_P1_More = 1'b0; $display(";A 6278");		//(= P2_P2_P1_More    0b0)) ;6278
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 6279");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b11101011)) ;6279
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 6280");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;6280
                                        if ((P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 6282");		//(= (bool-to-bv (bv-gt P2_P2_P1_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;6282
                                            P2_P2_P1_PhyAddrPointer = ((P2_P2_P1_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 6284");		//(= P2_P2_P1_PhyAddrPointer    (bv-sub (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P2_P2_P1_InstQueue 0 )))) ;6284
                                            P2_P2_P1_InstAddrPointer = P2_P2_P1_PhyAddrPointer; $display(";A 6285");		//(= P2_P2_P1_InstAddrPointer    P2_P2_P1_PhyAddrPointer )) ;6285
                                        end
                                        else begin
                                            $display(";A 6283");		//(= (bool-to-bv (bv-gt P2_P2_P1_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;6283
                                            P2_P2_P1_PhyAddrPointer = ((P2_P2_P1_InstAddrPointer + 32'b00000000000000000000000000000010) + P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 6286");		//(= P2_P2_P1_PhyAddrPointer    (bv-add (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000010) P2_P2_P1_InstQueue 0 ))) ;6286
                                            P2_P2_P1_InstAddrPointer = P2_P2_P1_PhyAddrPointer; $display(";A 6287");		//(= P2_P2_P1_InstAddrPointer    P2_P2_P1_PhyAddrPointer )) ;6287
                                        end
                                        P2_P2_P1_Flush = 1'b1; $display(";A 6288");		//(= P2_P2_P1_Flush    0b1)) ;6288
                                        P2_P2_P1_More = 1'b0; $display(";A 6289");		//(= P2_P2_P1_More    0b0)) ;6289
                                    end
                                    else begin
                                        $display(";A 6281");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;6281
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6290");		//(= P2_P2_P1_Flush    0b0)) ;6290
                                        P2_P2_P1_More = 1'b1; $display(";A 6291");		//(= P2_P2_P1_More    0b1)) ;6291
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 6292");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b11101001)) ;6292
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 6293");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;6293
                                        P2_P2_P1_PhyAddrPointer = ((P2_P2_P1_InstAddrPointer + 32'b00000000000000000000000000000101) + P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 6295");		//(= P2_P2_P1_PhyAddrPointer    (bv-add (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000101) P2_P2_P1_InstQueue 0 ))) ;6295
                                        P2_P2_P1_InstAddrPointer = P2_P2_P1_PhyAddrPointer; $display(";A 6296");		//(= P2_P2_P1_InstAddrPointer    P2_P2_P1_PhyAddrPointer )) ;6296
                                        P2_P2_P1_Flush = 1'b1; $display(";A 6297");		//(= P2_P2_P1_Flush    0b1)) ;6297
                                        P2_P2_P1_More = 1'b0; $display(";A 6298");		//(= P2_P2_P1_More    0b0)) ;6298
                                    end
                                    else begin
                                        $display(";A 6294");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;6294
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6299");		//(= P2_P2_P1_Flush    0b0)) ;6299
                                        P2_P2_P1_More = 1'b1; $display(";A 6300");		//(= P2_P2_P1_More    0b1)) ;6300
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 6301");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b11101010)) ;6301
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6302");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6302
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6303");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6303
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6304");		//(= P2_P2_P1_Flush    0b0)) ;6304
                                    P2_P2_P1_More = 1'b0; $display(";A 6305");		//(= P2_P2_P1_More    0b0)) ;6305
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 6306");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b10110000)) ;6306
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6307");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6307
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6308");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6308
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6309");		//(= P2_P2_P1_Flush    0b0)) ;6309
                                    P2_P2_P1_More = 1'b0; $display(";A 6310");		//(= P2_P2_P1_More    0b0)) ;6310
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 6311");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b10111000)) ;6311
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 6312");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;6312
                                        P2_P2_P1_EAX <= #1 ((((P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 6314");		//(= P2_P2_P1_EAX    (bv-add (bv-add (bv-add (bv-mul P2_P2_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P2_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P2_P1_InstQueue 0  0b00000000000000000000000100000000)) P2_P2_P1_InstQueue 0 ))) ;6314
                                        P2_P2_P1_More = 1'b0; $display(";A 6315");		//(= P2_P2_P1_More    0b0)) ;6315
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6316");		//(= P2_P2_P1_Flush    0b0)) ;6316
                                        P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 6317");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;6317
                                        P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 6318");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;6318
                                    end
                                    else begin
                                        $display(";A 6313");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;6313
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6319");		//(= P2_P2_P1_Flush    0b0)) ;6319
                                        P2_P2_P1_More = 1'b1; $display(";A 6320");		//(= P2_P2_P1_More    0b1)) ;6320
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 6321");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b10111011)) ;6321
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 6322");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;6322
                                        P2_P2_P1_EBX <= #1 ((((P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P2_P1_InstQueue[((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 6324");		//(= P2_P2_P1_EBX    (bv-add (bv-add (bv-add (bv-mul P2_P2_P1_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P2_P1_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P2_P1_InstQueue 0  0b00000000000000000000000100000000)) P2_P2_P1_InstQueue 0 ))) ;6324
                                        P2_P2_P1_More = 1'b0; $display(";A 6325");		//(= P2_P2_P1_More    0b0)) ;6325
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6326");		//(= P2_P2_P1_Flush    0b0)) ;6326
                                        P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 6327");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000101))) ;6327
                                        P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 6328");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;6328
                                    end
                                    else begin
                                        $display(";A 6323");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;6323
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6329");		//(= P2_P2_P1_Flush    0b0)) ;6329
                                        P2_P2_P1_More = 1'b1; $display(";A 6330");		//(= P2_P2_P1_More    0b1)) ;6330
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 6331");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b10001011)) ;6331
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6332");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6332
                                        if ((P2_P2_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 6334");		//(= (bool-to-bv (bv-slt P2_P2_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;6334
                                            P2_P2_P1_rEIP <= #1 (-P2_P2_P1_EBX); $display(";A 6336");		//(= P2_P2_P1_rEIP    (bv-neg P2_P2_P1_EBX ))) ;6336
                                        end
                                        else begin
                                            $display(";A 6335");		//(= (bool-to-bv (bv-slt P2_P2_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;6335
                                            P2_P2_P1_rEIP <= #1 P2_P2_P1_EBX; $display(";A 6337");		//(= P2_P2_P1_rEIP    P2_P2_P1_EBX )) ;6337
                                        end
                                        P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6338");		//(= P2_P2_P1_RequestPending    0b1)) ;6338
                                        P2_P2_P1_ReadRequest <= #1 1'b1; $display(";A 6339");		//(= P2_P2_P1_ReadRequest    0b1)) ;6339
                                        P2_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 6340");		//(= P2_P2_P1_MemoryFetch    0b1)) ;6340
                                        P2_P2_P1_CodeFetch <= #1 1'b0; $display(";A 6341");		//(= P2_P2_P1_CodeFetch    0b0)) ;6341
                                        if ((P2_P2_P1_READY_n == 1'b0)) begin
                                            $display(";A 6342");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6342
                                            P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6344");		//(= P2_P2_P1_RequestPending    0b0)) ;6344
                                            P2_P2_P1_uWord = (P2_P2_P1_Datai % 32'b00000000000000001000000000000000); $display(";A 6345");		//(= P2_P2_P1_uWord    (bv-smod P2_P2_P1_Datai  0b00000000000000001000000000000000))) ;6345
                                            if ((P2_P2_P1_StateBS16 == 1'b1)) begin
                                                $display(";A 6346");		//(= (bv-comp P2_P2_P1_StateBS16  0b1)   0b1)) ;6346
                                                P2_P2_P1_lWord = (P2_P2_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 6348");		//(= P2_P2_P1_lWord    (bv-smod P2_P2_P1_Datai  0b00000000000000010000000000000000))) ;6348
                                            end
                                            else begin
                                                $display(";A 6347");		//(= (bv-comp P2_P2_P1_StateBS16  0b1)   0b0)) ;6347
                                                P2_P2_P1_rEIP <= #1 (P2_P2_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 6349");		//(= P2_P2_P1_rEIP    (bv-add P2_P2_P1_rEIP  0b00000000000000000000000000000010))) ;6349
                                                P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6350");		//(= P2_P2_P1_RequestPending    0b1)) ;6350
                                                if ((P2_P2_P1_READY_n == 1'b0)) begin
                                                    $display(";A 6351");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6351
                                                    P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6353");		//(= P2_P2_P1_RequestPending    0b0)) ;6353
                                                    P2_P2_P1_lWord = (P2_P2_P1_Datai % 32'b00000000000000010000000000000000); $display(";A 6354");		//(= P2_P2_P1_lWord    (bv-smod P2_P2_P1_Datai  0b00000000000000010000000000000000))) ;6354
                                                end
                                                else begin
                                                    $display(";A 6352");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6352
                                                end
                                            end
                                            if ((P2_P2_P1_READY_n == 1'b0)) begin
                                                $display(";A 6355");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6355
                                                P2_P2_P1_EAX <= #1 ((P2_P2_P1_uWord * 32'b00000000000000010000000000000000) + P2_P2_P1_lWord); $display(";A 6357");		//(= P2_P2_P1_EAX    (bv-add (bv-mul P2_P2_P1_uWord  0b00000000000000010000000000000000) P2_P2_P1_lWord ))) ;6357
                                                P2_P2_P1_More = 1'b0; $display(";A 6358");		//(= P2_P2_P1_More    0b0)) ;6358
                                                P2_P2_P1_Flush = 1'b0; $display(";A 6359");		//(= P2_P2_P1_Flush    0b0)) ;6359
                                                P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6360");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;6360
                                                P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6361");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6361
                                            end
                                            else begin
                                                $display(";A 6356");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6356
                                            end
                                        end
                                        else begin
                                            $display(";A 6343");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6343
                                        end
                                    end
                                    else begin
                                        $display(";A 6333");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6333
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6362");		//(= P2_P2_P1_Flush    0b0)) ;6362
                                        P2_P2_P1_More = 1'b1; $display(";A 6363");		//(= P2_P2_P1_More    0b1)) ;6363
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 6364");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b10001001)) ;6364
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6365");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6365
                                        if ((P2_P2_P1_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 6367");		//(= (bool-to-bv (bv-slt P2_P2_P1_EBX  0b00000000000000000000000000000000))   0b1)) ;6367
                                            P2_P2_P1_rEIP <= #1 P2_P2_P1_EBX; $display(";A 6369");		//(= P2_P2_P1_rEIP    P2_P2_P1_EBX )) ;6369
                                        end
                                        else begin
                                            $display(";A 6368");		//(= (bool-to-bv (bv-slt P2_P2_P1_EBX  0b00000000000000000000000000000000))   0b0)) ;6368
                                            P2_P2_P1_rEIP <= #1 P2_P2_P1_EBX; $display(";A 6370");		//(= P2_P2_P1_rEIP    P2_P2_P1_EBX )) ;6370
                                        end
                                        P2_P2_P1_lWord = (P2_P2_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 6371");		//(= P2_P2_P1_lWord    (bv-smod P2_P2_P1_EAX  0b00000000000000010000000000000000))) ;6371
                                        P2_P2_P1_uWord = ((P2_P2_P1_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 6372");		//(= P2_P2_P1_uWord    (bv-smod (bv-sdiv P2_P2_P1_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;6372
                                        P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6373");		//(= P2_P2_P1_RequestPending    0b1)) ;6373
                                        P2_P2_P1_ReadRequest <= #1 1'b0; $display(";A 6374");		//(= P2_P2_P1_ReadRequest    0b0)) ;6374
                                        P2_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 6375");		//(= P2_P2_P1_MemoryFetch    0b1)) ;6375
                                        P2_P2_P1_CodeFetch <= #1 1'b0; $display(";A 6376");		//(= P2_P2_P1_CodeFetch    0b0)) ;6376
                                        if (((P2_P2_P1_State == 32'b00000000000000000000000000000010) | (P2_P2_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 6377");		//(= (bv-or (bv-comp P2_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P1_State  0b00000000000000000000000000000100))   0b1)) ;6377
                                            P2_P2_P1_Datao <= #1 ((P2_P2_P1_uWord * 32'b00000000000000010000000000000000) + P2_P2_P1_lWord); $display(";A 6379");		//(= P2_P2_P1_Datao    (bv-add (bv-mul P2_P2_P1_uWord  0b00000000000000010000000000000000) P2_P2_P1_lWord ))) ;6379
                                            if ((P2_P2_P1_READY_n == 1'b0)) begin
                                                $display(";A 6380");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6380
                                                P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6382");		//(= P2_P2_P1_RequestPending    0b0)) ;6382
                                                if ((P2_P2_P1_StateBS16 == 1'b0)) begin
                                                    $display(";A 6383");		//(= (bv-comp P2_P2_P1_StateBS16  0b0)   0b1)) ;6383
                                                    P2_P2_P1_rEIP <= #1 (P2_P2_P1_rEIP + 32'sb00000000000000000000000000000010); $display(";A 6385");		//(= P2_P2_P1_rEIP    (bv-add P2_P2_P1_rEIP  0b00000000000000000000000000000010))) ;6385
                                                    P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6386");		//(= P2_P2_P1_RequestPending    0b1)) ;6386
                                                    P2_P2_P1_ReadRequest <= #1 1'b0; $display(";A 6387");		//(= P2_P2_P1_ReadRequest    0b0)) ;6387
                                                    P2_P2_P1_MemoryFetch <= #1 1'b1; $display(";A 6388");		//(= P2_P2_P1_MemoryFetch    0b1)) ;6388
                                                    P2_P2_P1_CodeFetch <= #1 1'b0; $display(";A 6389");		//(= P2_P2_P1_CodeFetch    0b0)) ;6389
                                                    P2_P2_P1_State2 = 4'sb0110; $display(";A 6390");		//(= P2_P2_P1_State2    0b0110)) ;6390
                                                end
                                                else begin
                                                    $display(";A 6384");		//(= (bv-comp P2_P2_P1_StateBS16  0b0)   0b0)) ;6384
                                                end
                                                P2_P2_P1_More = 1'b0; $display(";A 6391");		//(= P2_P2_P1_More    0b0)) ;6391
                                                P2_P2_P1_Flush = 1'b0; $display(";A 6392");		//(= P2_P2_P1_Flush    0b0)) ;6392
                                                P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6393");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;6393
                                                P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6394");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6394
                                            end
                                            else begin
                                                $display(";A 6381");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6381
                                            end
                                        end
                                        else begin
                                            $display(";A 6378");		//(= (bv-or (bv-comp P2_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P1_State  0b00000000000000000000000000000100))   0b0)) ;6378
                                        end
                                    end
                                    else begin
                                        $display(";A 6366");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6366
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6395");		//(= P2_P2_P1_Flush    0b0)) ;6395
                                        P2_P2_P1_More = 1'b1; $display(";A 6396");		//(= P2_P2_P1_More    0b1)) ;6396
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 6397");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b11100100)) ;6397
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6398");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6398
                                        P2_P2_P1_rEIP <= #1 (P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 6400");		//(= P2_P2_P1_rEIP    (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;6400
                                        P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6401");		//(= P2_P2_P1_RequestPending    0b1)) ;6401
                                        P2_P2_P1_ReadRequest <= #1 1'b1; $display(";A 6402");		//(= P2_P2_P1_ReadRequest    0b1)) ;6402
                                        P2_P2_P1_MemoryFetch <= #1 1'b0; $display(";A 6403");		//(= P2_P2_P1_MemoryFetch    0b0)) ;6403
                                        P2_P2_P1_CodeFetch <= #1 1'b0; $display(";A 6404");		//(= P2_P2_P1_CodeFetch    0b0)) ;6404
                                        if ((P2_P2_P1_READY_n == 1'b0)) begin
                                            $display(";A 6405");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6405
                                            P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6407");		//(= P2_P2_P1_RequestPending    0b0)) ;6407
                                            P2_P2_P1_EAX <= #1 P2_P2_P1_Datai; $display(";A 6408");		//(= P2_P2_P1_EAX    P2_P2_P1_Datai )) ;6408
                                            P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6409");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;6409
                                            P2_P2_P1_InstQueueRd_Addr = (P2_P2_P1_InstQueueRd_Addr + 5'b00010); $display(";A 6410");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-add P2_P2_P1_InstQueueRd_Addr  0b00010))) ;6410
                                            P2_P2_P1_Flush = 1'b0; $display(";A 6411");		//(= P2_P2_P1_Flush    0b0)) ;6411
                                            P2_P2_P1_More = 1'b0; $display(";A 6412");		//(= P2_P2_P1_More    0b0)) ;6412
                                        end
                                        else begin
                                            $display(";A 6406");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6406
                                        end
                                    end
                                    else begin
                                        $display(";A 6399");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6399
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6413");		//(= P2_P2_P1_Flush    0b0)) ;6413
                                        P2_P2_P1_More = 1'b1; $display(";A 6414");		//(= P2_P2_P1_More    0b1)) ;6414
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 6415");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b11100110)) ;6415
                                    if (((P2_P2_P1_InstQueueWr_Addr - P2_P2_P1_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6416");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6416
                                        P2_P2_P1_rEIP <= #1 (P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 6418");		//(= P2_P2_P1_rEIP    (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;6418
                                        P2_P2_P1_RequestPending <= #1 1'b1; $display(";A 6419");		//(= P2_P2_P1_RequestPending    0b1)) ;6419
                                        P2_P2_P1_ReadRequest <= #1 1'b0; $display(";A 6420");		//(= P2_P2_P1_ReadRequest    0b0)) ;6420
                                        P2_P2_P1_MemoryFetch <= #1 1'b0; $display(";A 6421");		//(= P2_P2_P1_MemoryFetch    0b0)) ;6421
                                        P2_P2_P1_CodeFetch <= #1 1'b0; $display(";A 6422");		//(= P2_P2_P1_CodeFetch    0b0)) ;6422
                                        if (((P2_P2_P1_State == 32'b00000000000000000000000000000010) | (P2_P2_P1_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 6423");		//(= (bv-or (bv-comp P2_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P1_State  0b00000000000000000000000000000100))   0b1)) ;6423
                                            P2_P2_P1_fWord = (P2_P2_P1_EAX % 32'b00000000000000010000000000000000); $display(";A 6425");		//(= P2_P2_P1_fWord    (bv-smod P2_P2_P1_EAX  0b00000000000000010000000000000000))) ;6425
                                            P2_P2_P1_Datao <= #1 P2_P2_P1_fWord; $display(";A 6426");		//(= P2_P2_P1_Datao    P2_P2_P1_fWord )) ;6426
                                            if ((P2_P2_P1_READY_n == 1'b0)) begin
                                                $display(";A 6427");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6427
                                                P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6429");		//(= P2_P2_P1_RequestPending    0b0)) ;6429
                                                P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6430");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;6430
                                                P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6431");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6431
                                                P2_P2_P1_Flush = 1'b0; $display(";A 6432");		//(= P2_P2_P1_Flush    0b0)) ;6432
                                                P2_P2_P1_More = 1'b0; $display(";A 6433");		//(= P2_P2_P1_More    0b0)) ;6433
                                            end
                                            else begin
                                                $display(";A 6428");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6428
                                            end
                                        end
                                        else begin
                                            $display(";A 6424");		//(= (bv-or (bv-comp P2_P2_P1_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P1_State  0b00000000000000000000000000000100))   0b0)) ;6424
                                        end
                                    end
                                    else begin
                                        $display(";A 6417");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P1_InstQueueWr_Addr  P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6417
                                        P2_P2_P1_Flush = 1'b0; $display(";A 6434");		//(= P2_P2_P1_Flush    0b0)) ;6434
                                        P2_P2_P1_More = 1'b1; $display(";A 6435");		//(= P2_P2_P1_More    0b1)) ;6435
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 6436");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b00000100)) ;6436
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6437");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6437
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6438");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6438
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6439");		//(= P2_P2_P1_Flush    0b0)) ;6439
                                    P2_P2_P1_More = 1'b0; $display(";A 6440");		//(= P2_P2_P1_More    0b0)) ;6440
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 6441");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b00000101)) ;6441
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6442");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6442
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6443");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6443
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6444");		//(= P2_P2_P1_Flush    0b0)) ;6444
                                    P2_P2_P1_More = 1'b0; $display(";A 6445");		//(= P2_P2_P1_More    0b0)) ;6445
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 6446");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b11010000)) ;6446
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6447");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;6447
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6448");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6448
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6449");		//(= P2_P2_P1_Flush    0b0)) ;6449
                                    P2_P2_P1_More = 1'b0; $display(";A 6450");		//(= P2_P2_P1_More    0b0)) ;6450
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 6451");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b11000000)) ;6451
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6452");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000010))) ;6452
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6453");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6453
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6454");		//(= P2_P2_P1_Flush    0b0)) ;6454
                                    P2_P2_P1_More = 1'b0; $display(";A 6455");		//(= P2_P2_P1_More    0b0)) ;6455
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 6456");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b01000000)) ;6456
                                    P2_P2_P1_EAX <= #1 (P2_P2_P1_EAX + 32'sb00000000000000000000000000000001); $display(";A 6457");		//(= P2_P2_P1_EAX    (bv-add P2_P2_P1_EAX  0b00000000000000000000000000000001))) ;6457
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6458");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6458
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6459");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6459
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6460");		//(= P2_P2_P1_Flush    0b0)) ;6460
                                    P2_P2_P1_More = 1'b0; $display(";A 6461");		//(= P2_P2_P1_More    0b0)) ;6461
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 6462");		//(= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr )   0b01000011)) ;6462
                                    P2_P2_P1_EBX <= #1 (P2_P2_P1_EBX + 32'sb00000000000000000000000000000001); $display(";A 6463");		//(= P2_P2_P1_EBX    (bv-add P2_P2_P1_EBX  0b00000000000000000000000000000001))) ;6463
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6464");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6464
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6465");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6465
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6466");		//(= P2_P2_P1_Flush    0b0)) ;6466
                                    P2_P2_P1_More = 1'b0; $display(";A 6467");		//(= P2_P2_P1_More    0b0)) ;6467
                                end
                            default:
                                begin
                                    $display(";A 6468");		//(= (and (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b10010000) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b01100110) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b11101011) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b11101001) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b11101010) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b10110000) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b10111000) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b10111011) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b10001011) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b10001001) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b11100100) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b11100110) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b00000100) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b00000101) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b11010000) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b11000000) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b01000000) (/= ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ) 0b01000011))   true)) ;6468
                                    P2_P2_P1_InstAddrPointer = (P2_P2_P1_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6469");		//(= P2_P2_P1_InstAddrPointer    (bv-add P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000001))) ;6469
                                    P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6470");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6470
                                    P2_P2_P1_Flush = 1'b0; $display(";A 6471");		//(= P2_P2_P1_Flush    0b0)) ;6471
                                    P2_P2_P1_More = 1'b0; $display(";A 6472");		//(= P2_P2_P1_More    0b0)) ;6472
                                end
                        endcase
                        if (((~(P2_P2_P1_InstQueueRd_Addr < P2_P2_P1_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P2_P2_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P2_P2_P1_Flush) | P2_P2_P1_More))) begin
                            $display(";A 6473");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P2_P1_InstQueueRd_Addr  P2_P2_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P2_P1_Flush ) P2_P2_P1_More ))   0b1)) ;6473
                            P2_P2_P1_State2 = 4'sb0111; $display(";A 6475");		//(= P2_P2_P1_State2    0b0111)) ;6475
                        end
                        else begin
                            $display(";A 6474");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P2_P1_InstQueueRd_Addr  P2_P2_P1_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P2_P1_Flush ) P2_P2_P1_More ))   0b0)) ;6474
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 6476");		//(= P2_P2_P1_State2    0b0110)) ;6476
                        P2_P2_P1_Datao <= #1 ((P2_P2_P1_uWord * 32'b00000000000000010000000000000000) + P2_P2_P1_lWord); $display(";A 6477");		//(= P2_P2_P1_Datao    (bv-add (bv-mul P2_P2_P1_uWord  0b00000000000000010000000000000000) P2_P2_P1_lWord ))) ;6477
                        if ((P2_P2_P1_READY_n == 1'b0)) begin
                            $display(";A 6478");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b1)) ;6478
                            P2_P2_P1_RequestPending <= #1 1'b0; $display(";A 6480");		//(= P2_P2_P1_RequestPending    0b0)) ;6480
                            P2_P2_P1_State2 = 4'sb0101; $display(";A 6481");		//(= P2_P2_P1_State2    0b0101)) ;6481
                        end
                        else begin
                            $display(";A 6479");		//(= (bv-comp P2_P2_P1_READY_n  0b0)   0b0)) ;6479
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 6482");		//(= P2_P2_P1_State2    0b0111)) ;6482
                        if (P2_P2_P1_Flush) begin
                            $display(";A 6483");		//(= P2_P2_P1_Flush    0b1)) ;6483
                            P2_P2_P1_InstQueueRd_Addr = 5'sb00001; $display(";A 6485");		//(= P2_P2_P1_InstQueueRd_Addr    0b00001)) ;6485
                            P2_P2_P1_InstQueueWr_Addr = 5'sb00001; $display(";A 6486");		//(= P2_P2_P1_InstQueueWr_Addr    0b00001)) ;6486
                            if ((P2_P2_P1_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 6487");		//(= (bool-to-bv (bv-slt P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;6487
                                P2_P2_P1_fWord = (-P2_P2_P1_InstAddrPointer); $display(";A 6489");		//(= P2_P2_P1_fWord    (bv-neg P2_P2_P1_InstAddrPointer ))) ;6489
                            end
                            else begin
                                $display(";A 6488");		//(= (bool-to-bv (bv-slt P2_P2_P1_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;6488
                                P2_P2_P1_fWord = P2_P2_P1_InstAddrPointer; $display(";A 6490");		//(= P2_P2_P1_fWord    P2_P2_P1_InstAddrPointer )) ;6490
                            end
                            if (((P2_P2_P1_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 6491");		//(= (bv-comp (bv-smod P2_P2_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;6491
                                P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + (P2_P2_P1_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 6493");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  (bv-smod P2_P2_P1_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;6493
                            end
                            else begin
                                $display(";A 6492");		//(= (bv-comp (bv-smod P2_P2_P1_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;6492
                            end
                        end
                        else begin
                            $display(";A 6484");		//(= P2_P2_P1_Flush    0b0)) ;6484
                        end
                        if (((32'b00000000000000000000000000001111 - P2_P2_P1_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 6494");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;6494
                            P2_P2_P1_State2 = 4'sb1000; $display(";A 6496");		//(= P2_P2_P1_State2    0b1000)) ;6496
                            P2_P2_P1_InstQueueWr_Addr = 5'sb00000; $display(";A 6497");		//(= P2_P2_P1_InstQueueWr_Addr    0b00000)) ;6497
                        end
                        else begin
                            $display(";A 6495");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P1_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;6495
                            P2_P2_P1_State2 = 4'sb1001; $display(";A 6498");		//(= P2_P2_P1_State2    0b1001)) ;6498
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 6499");		//(= P2_P2_P1_State2    0b1000)) ;6499
                        if ((P2_P2_P1_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 6500");		//(= (bool-to-bv (bv-le P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;6500
                            P2_P2_P1_InstQueue[P2_P2_P1_InstQueueWr_Addr] = P2_P2_P1_InstQueue[P2_P2_P1_InstQueueRd_Addr]; $display(";A 6502");		//(= P2_P2_P1_InstQueue    ( P2_P2_P1_InstQueue P2_P2_P1_InstQueueRd_Addr ))) ;6502
                            P2_P2_P1_InstQueueRd_Addr = ((P2_P2_P1_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6503");		//(= P2_P2_P1_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6503
                            P2_P2_P1_InstQueueWr_Addr = ((P2_P2_P1_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6504");		//(= P2_P2_P1_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P1_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6504
                            P2_P2_P1_State2 = 4'sb1000; $display(";A 6505");		//(= P2_P2_P1_State2    0b1000)) ;6505
                        end
                        else begin
                            $display(";A 6501");		//(= (bool-to-bv (bv-le P2_P2_P1_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;6501
                            P2_P2_P1_InstQueueRd_Addr = 5'sb00000; $display(";A 6506");		//(= P2_P2_P1_InstQueueRd_Addr    0b00000)) ;6506
                            P2_P2_P1_State2 = 4'sb1001; $display(";A 6507");		//(= P2_P2_P1_State2    0b1001)) ;6507
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 6508");		//(= P2_P2_P1_State2    0b1001)) ;6508
                        P2_P2_P1_rEIP <= #1 P2_P2_P1_PhyAddrPointer; $display(";A 6509");		//(= P2_P2_P1_rEIP    P2_P2_P1_PhyAddrPointer )) ;6509
                        P2_P2_P1_State2 = 4'sb0001; $display(";A 6510");		//(= P2_P2_P1_State2    0b0001)) ;6510
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:9945
    always @(posedge P2_P2_P1_RESET or posedge P2_P2_P1_CLOCK) begin
        if ((P2_P2_P1_RESET == 1'b1)) begin
            $display(";A 6511");		//(= (bv-comp P2_P2_P1_RESET  0b1)   0b1)) ;6511
            P2_P2_P1_ByteEnable <= #1 4'b0000; $display(";A 6513");		//(= P2_P2_P1_ByteEnable    0b0000)) ;6513
            P2_P2_P1_NonAligned <= #1 1'b0; $display(";A 6514");		//(= P2_P2_P1_NonAligned    0b0)) ;6514
        end
        else begin
            $display(";A 6512");		//(= (bv-comp P2_P2_P1_RESET  0b1)   0b0)) ;6512
            case (P2_P2_P1_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 6515");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000000)) ;6515
                        case ((P2_P2_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 6516");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;6516
                                    P2_P2_P1_ByteEnable <= #1 4'b1110; $display(";A 6517");		//(= P2_P2_P1_ByteEnable    0b1110)) ;6517
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 6518");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;6518
                                    P2_P2_P1_ByteEnable <= #1 4'b1101; $display(";A 6519");		//(= P2_P2_P1_ByteEnable    0b1101)) ;6519
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 6520");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;6520
                                    P2_P2_P1_ByteEnable <= #1 4'b1011; $display(";A 6521");		//(= P2_P2_P1_ByteEnable    0b1011)) ;6521
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 6522");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;6522
                                    P2_P2_P1_ByteEnable <= #1 4'b0111; $display(";A 6523");		//(= P2_P2_P1_ByteEnable    0b0111)) ;6523
                                end
                            default:
                                begin
                                    $display(";A 6524");		//(= (and (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;6524
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 6525");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000001)) ;6525
                        case ((P2_P2_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 6526");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;6526
                                    P2_P2_P1_ByteEnable <= #1 4'b1100; $display(";A 6527");		//(= P2_P2_P1_ByteEnable    0b1100)) ;6527
                                    P2_P2_P1_NonAligned <= #1 1'b0; $display(";A 6528");		//(= P2_P2_P1_NonAligned    0b0)) ;6528
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 6529");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;6529
                                    P2_P2_P1_ByteEnable <= #1 4'b1001; $display(";A 6530");		//(= P2_P2_P1_ByteEnable    0b1001)) ;6530
                                    P2_P2_P1_NonAligned <= #1 1'b0; $display(";A 6531");		//(= P2_P2_P1_NonAligned    0b0)) ;6531
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 6532");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;6532
                                    P2_P2_P1_ByteEnable <= #1 4'b0011; $display(";A 6533");		//(= P2_P2_P1_ByteEnable    0b0011)) ;6533
                                    P2_P2_P1_NonAligned <= #1 1'b0; $display(";A 6534");		//(= P2_P2_P1_NonAligned    0b0)) ;6534
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 6535");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;6535
                                    P2_P2_P1_ByteEnable <= #1 4'b0111; $display(";A 6536");		//(= P2_P2_P1_ByteEnable    0b0111)) ;6536
                                    P2_P2_P1_NonAligned <= #1 1'b1; $display(";A 6537");		//(= P2_P2_P1_NonAligned    0b1)) ;6537
                                end
                            default:
                                begin
                                    $display(";A 6538");		//(= (and (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;6538
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 6539");		//(= P2_P2_P1_DataWidth    0b00000000000000000000000000000010)) ;6539
                        case ((P2_P2_P1_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 6540");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;6540
                                    P2_P2_P1_ByteEnable <= #1 4'b0000; $display(";A 6541");		//(= P2_P2_P1_ByteEnable    0b0000)) ;6541
                                    P2_P2_P1_NonAligned <= #1 1'b0; $display(";A 6542");		//(= P2_P2_P1_NonAligned    0b0)) ;6542
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 6543");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;6543
                                    P2_P2_P1_ByteEnable <= #1 4'b0001; $display(";A 6544");		//(= P2_P2_P1_ByteEnable    0b0001)) ;6544
                                    P2_P2_P1_NonAligned <= #1 1'b1; $display(";A 6545");		//(= P2_P2_P1_NonAligned    0b1)) ;6545
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 6546");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;6546
                                    P2_P2_P1_NonAligned <= #1 1'b1; $display(";A 6547");		//(= P2_P2_P1_NonAligned    0b1)) ;6547
                                    P2_P2_P1_ByteEnable <= #1 4'b0011; $display(";A 6548");		//(= P2_P2_P1_ByteEnable    0b0011)) ;6548
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 6549");		//(= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;6549
                                    P2_P2_P1_NonAligned <= #1 1'b1; $display(";A 6550");		//(= P2_P2_P1_NonAligned    0b1)) ;6550
                                    P2_P2_P1_ByteEnable <= #1 4'b0111; $display(";A 6551");		//(= P2_P2_P1_ByteEnable    0b0111)) ;6551
                                end
                            default:
                                begin
                                    $display(";A 6552");		//(= (and (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P1_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;6552
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 6553");		//(= (and (/= P2_P2_P1_DataWidth  0b00000000000000000000000000000000) (/= P2_P2_P1_DataWidth  0b00000000000000000000000000000001) (/= P2_P2_P1_DataWidth  0b00000000000000000000000000000010))   true)) ;6553
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:10133
    always @(posedge P2_P2_P2_RESET or posedge P2_P2_P2_CLOCK) begin
        if ((P2_P2_P2_RESET == 1'b1)) begin
            $display(";A 6554");		//(= (bv-comp P2_P2_P2_RESET  0b1)   0b1)) ;6554
            P2_P2_P2_BE_n <= #1 4'b0000; $display(";A 6556");		//(= P2_P2_P2_BE_n    0b0000)) ;6556
            P2_P2_P2_Address <= #1 30'sb000000000000000000000000000000; $display(";A 6557");		//(= P2_P2_P2_Address    0b000000000000000000000000000000)) ;6557
            P2_P2_P2_W_R_n <= #1 1'b0; $display(";A 6558");		//(= P2_P2_P2_W_R_n    0b0)) ;6558
            P2_P2_P2_D_C_n <= #1 1'b0; $display(";A 6559");		//(= P2_P2_P2_D_C_n    0b0)) ;6559
            P2_P2_P2_M_IO_n <= #1 1'b0; $display(";A 6560");		//(= P2_P2_P2_M_IO_n    0b0)) ;6560
            P2_P2_P2_ADS_n <= #1 1'b0; $display(";A 6561");		//(= P2_P2_P2_ADS_n    0b0)) ;6561
            P2_P2_P2_State <= #1 3'sb000; $display(";A 6562");		//(= P2_P2_P2_State    0b000)) ;6562
            P2_P2_P2_StateNA <= #1 1'b0; $display(";A 6563");		//(= P2_P2_P2_StateNA    0b0)) ;6563
            P2_P2_P2_StateBS16 <= #1 1'b0; $display(";A 6564");		//(= P2_P2_P2_StateBS16    0b0)) ;6564
            P2_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 6565");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000000)) ;6565
        end
        else begin
            $display(";A 6555");		//(= (bv-comp P2_P2_P2_RESET  0b1)   0b0)) ;6555
            case (P2_P2_P2_State)
                3'b000 :
                    begin
                        $display(";A 6566");		//(= P2_P2_P2_State    0b000)) ;6566
                        P2_P2_P2_D_C_n <= #1 1'b1; $display(";A 6567");		//(= P2_P2_P2_D_C_n    0b1)) ;6567
                        P2_P2_P2_ADS_n <= #1 1'b1; $display(";A 6568");		//(= P2_P2_P2_ADS_n    0b1)) ;6568
                        P2_P2_P2_State <= #1 3'sb001; $display(";A 6569");		//(= P2_P2_P2_State    0b001)) ;6569
                        P2_P2_P2_StateNA <= #1 1'b1; $display(";A 6570");		//(= P2_P2_P2_StateNA    0b1)) ;6570
                        P2_P2_P2_StateBS16 <= #1 1'b1; $display(";A 6571");		//(= P2_P2_P2_StateBS16    0b1)) ;6571
                        P2_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 6572");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;6572
                        P2_P2_P2_State <= #1 3'sb001; $display(";A 6573");		//(= P2_P2_P2_State    0b001)) ;6573
                    end
                3'b001 :
                    begin
                        $display(";A 6574");		//(= P2_P2_P2_State    0b001)) ;6574
                        if ((P2_P2_P2_RequestPending == 1'b1)) begin
                            $display(";A 6575");		//(= (bv-comp P2_P2_P2_RequestPending  0b1)   0b1)) ;6575
                            P2_P2_P2_State <= #1 3'sb010; $display(";A 6577");		//(= P2_P2_P2_State    0b010)) ;6577
                        end
                        else begin
                            $display(";A 6576");		//(= (bv-comp P2_P2_P2_RequestPending  0b1)   0b0)) ;6576
                            if ((P2_P2_P2_HOLD == 1'b1)) begin
                                $display(";A 6578");		//(= (bv-comp P2_P2_P2_HOLD  0b1)   0b1)) ;6578
                                P2_P2_P2_State <= #1 3'sb101; $display(";A 6580");		//(= P2_P2_P2_State    0b101)) ;6580
                            end
                            else begin
                                $display(";A 6579");		//(= (bv-comp P2_P2_P2_HOLD  0b1)   0b0)) ;6579
                                P2_P2_P2_State <= #1 3'sb001; $display(";A 6581");		//(= P2_P2_P2_State    0b001)) ;6581
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 6582");		//(= P2_P2_P2_State    0b010)) ;6582
                        P2_P2_P2_Address <= #1 ((P2_P2_P2_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 6583");		//(= P2_P2_P2_Address    (bv-smod (bv-sdiv P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;6583
                        P2_P2_P2_BE_n <= #1 P2_P2_P2_ByteEnable; $display(";A 6584");		//(= P2_P2_P2_BE_n    P2_P2_P2_ByteEnable )) ;6584
                        P2_P2_P2_M_IO_n <= #1 P2_P2_P2_MemoryFetch; $display(";A 6585");		//(= P2_P2_P2_M_IO_n    P2_P2_P2_MemoryFetch )) ;6585
                        if ((P2_P2_P2_ReadRequest == 1'b1)) begin
                            $display(";A 6586");		//(= (bv-comp P2_P2_P2_ReadRequest  0b1)   0b1)) ;6586
                            P2_P2_P2_W_R_n <= #1 1'b0; $display(";A 6588");		//(= P2_P2_P2_W_R_n    0b0)) ;6588
                        end
                        else begin
                            $display(";A 6587");		//(= (bv-comp P2_P2_P2_ReadRequest  0b1)   0b0)) ;6587
                            P2_P2_P2_W_R_n <= #1 1'b1; $display(";A 6589");		//(= P2_P2_P2_W_R_n    0b1)) ;6589
                        end
                        if ((P2_P2_P2_CodeFetch == 1'b1)) begin
                            $display(";A 6590");		//(= (bv-comp P2_P2_P2_CodeFetch  0b1)   0b1)) ;6590
                            P2_P2_P2_D_C_n <= #1 1'b0; $display(";A 6592");		//(= P2_P2_P2_D_C_n    0b0)) ;6592
                        end
                        else begin
                            $display(";A 6591");		//(= (bv-comp P2_P2_P2_CodeFetch  0b1)   0b0)) ;6591
                            P2_P2_P2_D_C_n <= #1 1'b1; $display(";A 6593");		//(= P2_P2_P2_D_C_n    0b1)) ;6593
                        end
                        P2_P2_P2_ADS_n <= #1 1'b0; $display(";A 6594");		//(= P2_P2_P2_ADS_n    0b0)) ;6594
                        P2_P2_P2_State <= #1 3'sb011; $display(";A 6595");		//(= P2_P2_P2_State    0b011)) ;6595
                    end
                3'b011 :
                    begin
                        $display(";A 6596");		//(= P2_P2_P2_State    0b011)) ;6596
                        if ((((P2_P2_P2_READY_n == 1'b0) & (P2_P2_P2_HOLD == 1'b0)) & (P2_P2_P2_RequestPending == 1'b1))) begin
                            $display(";A 6597");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b1))   0b1)) ;6597
                            P2_P2_P2_State <= #1 3'sb010; $display(";A 6599");		//(= P2_P2_P2_State    0b010)) ;6599
                        end
                        else begin
                            $display(";A 6598");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b1))   0b0)) ;6598
                            if (((P2_P2_P2_READY_n == 1'b1) & (P2_P2_P2_NA_n == 1'b1))) begin
                                $display(";A 6600");		//(= (bv-and (bv-comp P2_P2_P2_READY_n  0b1) (bv-comp P2_P2_P2_NA_n  0b1))   0b1)) ;6600
                            end
                            else begin
                                $display(";A 6601");		//(= (bv-and (bv-comp P2_P2_P2_READY_n  0b1) (bv-comp P2_P2_P2_NA_n  0b1))   0b0)) ;6601
                                if ((((P2_P2_P2_RequestPending == 1'b1) | (P2_P2_P2_HOLD == 1'b1)) & ((P2_P2_P2_READY_n == 1'b1) & (P2_P2_P2_NA_n == 1'b0)))) begin
                                    $display(";A 6602");		//(= (bv-and (bv-or (bv-comp P2_P2_P2_RequestPending  0b1) (bv-comp P2_P2_P2_HOLD  0b1)) (bv-and (bv-comp P2_P2_P2_READY_n  0b1) (bv-comp P2_P2_P2_NA_n  0b0)))   0b1)) ;6602
                                    P2_P2_P2_State <= #1 3'sb111; $display(";A 6604");		//(= P2_P2_P2_State    0b111)) ;6604
                                end
                                else begin
                                    $display(";A 6603");		//(= (bv-and (bv-or (bv-comp P2_P2_P2_RequestPending  0b1) (bv-comp P2_P2_P2_HOLD  0b1)) (bv-and (bv-comp P2_P2_P2_READY_n  0b1) (bv-comp P2_P2_P2_NA_n  0b0)))   0b0)) ;6603
                                    if (((((P2_P2_P2_RequestPending == 1'b1) & (P2_P2_P2_HOLD == 1'b0)) & (P2_P2_P2_READY_n == 1'b1)) & (P2_P2_P2_NA_n == 1'b0))) begin
                                        $display(";A 6605");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P2_P2_RequestPending  0b1) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_READY_n  0b1)) (bv-comp P2_P2_P2_NA_n  0b0))   0b1)) ;6605
                                        P2_P2_P2_State <= #1 3'sb110; $display(";A 6607");		//(= P2_P2_P2_State    0b110)) ;6607
                                    end
                                    else begin
                                        $display(";A 6606");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P2_P2_RequestPending  0b1) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_READY_n  0b1)) (bv-comp P2_P2_P2_NA_n  0b0))   0b0)) ;6606
                                        if ((((P2_P2_P2_RequestPending == 1'b0) & (P2_P2_P2_HOLD == 1'b0)) & (P2_P2_P2_READY_n == 1'b0))) begin
                                            $display(";A 6608");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_RequestPending  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_READY_n  0b0))   0b1)) ;6608
                                            P2_P2_P2_State <= #1 3'sb001; $display(";A 6610");		//(= P2_P2_P2_State    0b001)) ;6610
                                        end
                                        else begin
                                            $display(";A 6609");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_RequestPending  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_READY_n  0b0))   0b0)) ;6609
                                            if (((P2_P2_P2_HOLD == 1'b1) & (P2_P2_P2_READY_n == 1'b1))) begin
                                                $display(";A 6611");		//(= (bv-and (bv-comp P2_P2_P2_HOLD  0b1) (bv-comp P2_P2_P2_READY_n  0b1))   0b1)) ;6611
                                                P2_P2_P2_State <= #1 3'sb101; $display(";A 6613");		//(= P2_P2_P2_State    0b101)) ;6613
                                            end
                                            else begin
                                                $display(";A 6612");		//(= (bv-and (bv-comp P2_P2_P2_HOLD  0b1) (bv-comp P2_P2_P2_READY_n  0b1))   0b0)) ;6612
                                                P2_P2_P2_State <= #1 3'sb011; $display(";A 6614");		//(= P2_P2_P2_State    0b011)) ;6614
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P2_P2_P2_StateBS16 <= #1 P2_P2_P2_BS16_n; $display(";A 6615");		//(= P2_P2_P2_StateBS16    P2_P2_P2_BS16_n )) ;6615
                        if ((P2_P2_P2_BS16_n == 1'b0)) begin
                            $display(";A 6616");		//(= (bv-comp P2_P2_P2_BS16_n  0b0)   0b1)) ;6616
                            P2_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 6618");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000001)) ;6618
                        end
                        else begin
                            $display(";A 6617");		//(= (bv-comp P2_P2_P2_BS16_n  0b0)   0b0)) ;6617
                            P2_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 6619");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;6619
                        end
                        P2_P2_P2_StateNA <= #1 P2_P2_P2_NA_n; $display(";A 6620");		//(= P2_P2_P2_StateNA    P2_P2_P2_NA_n )) ;6620
                        P2_P2_P2_ADS_n <= #1 1'b1; $display(";A 6621");		//(= P2_P2_P2_ADS_n    0b1)) ;6621
                    end
                3'b100 :
                    begin
                        $display(";A 6622");		//(= P2_P2_P2_State    0b100)) ;6622
                        if ((((P2_P2_P2_NA_n == 1'b0) & (P2_P2_P2_HOLD == 1'b0)) & (P2_P2_P2_RequestPending == 1'b1))) begin
                            $display(";A 6623");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_NA_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b1))   0b1)) ;6623
                            P2_P2_P2_State <= #1 3'sb110; $display(";A 6625");		//(= P2_P2_P2_State    0b110)) ;6625
                        end
                        else begin
                            $display(";A 6624");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_NA_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b1))   0b0)) ;6624
                            if (((P2_P2_P2_NA_n == 1'b0) & ((P2_P2_P2_HOLD == 1'b1) | (P2_P2_P2_RequestPending == 1'b0)))) begin
                                $display(";A 6626");		//(= (bv-and (bv-comp P2_P2_P2_NA_n  0b0) (bv-or (bv-comp P2_P2_P2_HOLD  0b1) (bv-comp P2_P2_P2_RequestPending  0b0)))   0b1)) ;6626
                                P2_P2_P2_State <= #1 3'sb111; $display(";A 6628");		//(= P2_P2_P2_State    0b111)) ;6628
                            end
                            else begin
                                $display(";A 6627");		//(= (bv-and (bv-comp P2_P2_P2_NA_n  0b0) (bv-or (bv-comp P2_P2_P2_HOLD  0b1) (bv-comp P2_P2_P2_RequestPending  0b0)))   0b0)) ;6627
                                if ((P2_P2_P2_NA_n == 1'b1)) begin
                                    $display(";A 6629");		//(= (bv-comp P2_P2_P2_NA_n  0b1)   0b1)) ;6629
                                    P2_P2_P2_State <= #1 3'sb011; $display(";A 6631");		//(= P2_P2_P2_State    0b011)) ;6631
                                end
                                else begin
                                    $display(";A 6630");		//(= (bv-comp P2_P2_P2_NA_n  0b1)   0b0)) ;6630
                                    P2_P2_P2_State <= #1 3'sb100; $display(";A 6632");		//(= P2_P2_P2_State    0b100)) ;6632
                                end
                            end
                        end
                        P2_P2_P2_StateBS16 <= #1 P2_P2_P2_BS16_n; $display(";A 6633");		//(= P2_P2_P2_StateBS16    P2_P2_P2_BS16_n )) ;6633
                        if ((P2_P2_P2_BS16_n == 1'b0)) begin
                            $display(";A 6634");		//(= (bv-comp P2_P2_P2_BS16_n  0b0)   0b1)) ;6634
                            P2_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 6636");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000001)) ;6636
                        end
                        else begin
                            $display(";A 6635");		//(= (bv-comp P2_P2_P2_BS16_n  0b0)   0b0)) ;6635
                            P2_P2_P2_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 6637");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;6637
                        end
                        P2_P2_P2_StateNA <= #1 P2_P2_P2_NA_n; $display(";A 6638");		//(= P2_P2_P2_StateNA    P2_P2_P2_NA_n )) ;6638
                        P2_P2_P2_ADS_n <= #1 1'b1; $display(";A 6639");		//(= P2_P2_P2_ADS_n    0b1)) ;6639
                    end
                3'b101 :
                    begin
                        $display(";A 6640");		//(= P2_P2_P2_State    0b101)) ;6640
                        if (((P2_P2_P2_HOLD == 1'b0) & (P2_P2_P2_RequestPending == 1'b1))) begin
                            $display(";A 6641");		//(= (bv-and (bv-comp P2_P2_P2_HOLD  0b0) (bv-comp P2_P2_P2_RequestPending  0b1))   0b1)) ;6641
                            P2_P2_P2_State <= #1 3'sb010; $display(";A 6643");		//(= P2_P2_P2_State    0b010)) ;6643
                        end
                        else begin
                            $display(";A 6642");		//(= (bv-and (bv-comp P2_P2_P2_HOLD  0b0) (bv-comp P2_P2_P2_RequestPending  0b1))   0b0)) ;6642
                            if (((P2_P2_P2_HOLD == 1'b0) & (P2_P2_P2_RequestPending == 1'b0))) begin
                                $display(";A 6644");		//(= (bv-and (bv-comp P2_P2_P2_HOLD  0b0) (bv-comp P2_P2_P2_RequestPending  0b0))   0b1)) ;6644
                                P2_P2_P2_State <= #1 3'sb001; $display(";A 6646");		//(= P2_P2_P2_State    0b001)) ;6646
                            end
                            else begin
                                $display(";A 6645");		//(= (bv-and (bv-comp P2_P2_P2_HOLD  0b0) (bv-comp P2_P2_P2_RequestPending  0b0))   0b0)) ;6645
                                P2_P2_P2_State <= #1 3'sb101; $display(";A 6647");		//(= P2_P2_P2_State    0b101)) ;6647
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 6648");		//(= P2_P2_P2_State    0b110)) ;6648
                        P2_P2_P2_Address <= #1 ((P2_P2_P2_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 6649");		//(= P2_P2_P2_Address    (bv-smod (bv-sdiv P2_P2_P2_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;6649
                        P2_P2_P2_BE_n <= #1 P2_P2_P2_ByteEnable; $display(";A 6650");		//(= P2_P2_P2_BE_n    P2_P2_P2_ByteEnable )) ;6650
                        P2_P2_P2_M_IO_n <= #1 P2_P2_P2_MemoryFetch; $display(";A 6651");		//(= P2_P2_P2_M_IO_n    P2_P2_P2_MemoryFetch )) ;6651
                        if ((P2_P2_P2_ReadRequest == 1'b1)) begin
                            $display(";A 6652");		//(= (bv-comp P2_P2_P2_ReadRequest  0b1)   0b1)) ;6652
                            P2_P2_P2_W_R_n <= #1 1'b0; $display(";A 6654");		//(= P2_P2_P2_W_R_n    0b0)) ;6654
                        end
                        else begin
                            $display(";A 6653");		//(= (bv-comp P2_P2_P2_ReadRequest  0b1)   0b0)) ;6653
                            P2_P2_P2_W_R_n <= #1 1'b1; $display(";A 6655");		//(= P2_P2_P2_W_R_n    0b1)) ;6655
                        end
                        if ((P2_P2_P2_CodeFetch == 1'b1)) begin
                            $display(";A 6656");		//(= (bv-comp P2_P2_P2_CodeFetch  0b1)   0b1)) ;6656
                            P2_P2_P2_D_C_n <= #1 1'b0; $display(";A 6658");		//(= P2_P2_P2_D_C_n    0b0)) ;6658
                        end
                        else begin
                            $display(";A 6657");		//(= (bv-comp P2_P2_P2_CodeFetch  0b1)   0b0)) ;6657
                            P2_P2_P2_D_C_n <= #1 1'b1; $display(";A 6659");		//(= P2_P2_P2_D_C_n    0b1)) ;6659
                        end
                        P2_P2_P2_ADS_n <= #1 1'b0; $display(";A 6660");		//(= P2_P2_P2_ADS_n    0b0)) ;6660
                        if ((P2_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 6661");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6661
                            P2_P2_P2_State <= #1 3'sb100; $display(";A 6663");		//(= P2_P2_P2_State    0b100)) ;6663
                        end
                        else begin
                            $display(";A 6662");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6662
                            P2_P2_P2_State <= #1 3'sb110; $display(";A 6664");		//(= P2_P2_P2_State    0b110)) ;6664
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 6665");		//(= P2_P2_P2_State    0b111)) ;6665
                        if ((((P2_P2_P2_READY_n == 1'b1) & (P2_P2_P2_RequestPending == 1'b1)) & (P2_P2_P2_HOLD == 1'b0))) begin
                            $display(";A 6666");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b1) (bv-comp P2_P2_P2_RequestPending  0b1)) (bv-comp P2_P2_P2_HOLD  0b0))   0b1)) ;6666
                            P2_P2_P2_State <= #1 3'sb110; $display(";A 6668");		//(= P2_P2_P2_State    0b110)) ;6668
                        end
                        else begin
                            $display(";A 6667");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b1) (bv-comp P2_P2_P2_RequestPending  0b1)) (bv-comp P2_P2_P2_HOLD  0b0))   0b0)) ;6667
                            if (((P2_P2_P2_READY_n == 1'b0) & (P2_P2_P2_HOLD == 1'b1))) begin
                                $display(";A 6669");		//(= (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b1))   0b1)) ;6669
                                P2_P2_P2_State <= #1 3'sb101; $display(";A 6671");		//(= P2_P2_P2_State    0b101)) ;6671
                            end
                            else begin
                                $display(";A 6670");		//(= (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b1))   0b0)) ;6670
                                if ((((P2_P2_P2_READY_n == 1'b0) & (P2_P2_P2_HOLD == 1'b0)) & (P2_P2_P2_RequestPending == 1'b1))) begin
                                    $display(";A 6672");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b1))   0b1)) ;6672
                                    P2_P2_P2_State <= #1 3'sb010; $display(";A 6674");		//(= P2_P2_P2_State    0b010)) ;6674
                                end
                                else begin
                                    $display(";A 6673");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b1))   0b0)) ;6673
                                    if ((((P2_P2_P2_READY_n == 1'b0) & (P2_P2_P2_HOLD == 1'b0)) & (P2_P2_P2_RequestPending == 1'b0))) begin
                                        $display(";A 6675");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b0))   0b1)) ;6675
                                        P2_P2_P2_State <= #1 3'sb001; $display(";A 6677");		//(= P2_P2_P2_State    0b001)) ;6677
                                    end
                                    else begin
                                        $display(";A 6676");		//(= (bv-and (bv-and (bv-comp P2_P2_P2_READY_n  0b0) (bv-comp P2_P2_P2_HOLD  0b0)) (bv-comp P2_P2_P2_RequestPending  0b0))   0b0)) ;6676
                                        P2_P2_P2_State <= #1 3'sb111; $display(";A 6678");		//(= P2_P2_P2_State    0b111)) ;6678
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:10277
    always @(posedge P2_P2_P2_RESET or posedge P2_P2_P2_CLOCK) begin
        if ((P2_P2_P2_RESET == 1'b1)) begin
            $display(";A 6679");		//(= (bv-comp P2_P2_P2_RESET  0b1)   0b1)) ;6679
            P2_P2_P2_State2 = 4'sb0000; $display(";A 6681");		//(= P2_P2_P2_State2    0b0000)) ;6681
            P2_P2_P2_InstQueue[0] = 8'b00000000; $display(";A 6682");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6682
            P2_P2_P2_InstQueue[1] = 8'b00000000; $display(";A 6683");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6683
            P2_P2_P2_InstQueue[2] = 8'b00000000; $display(";A 6684");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6684
            P2_P2_P2_InstQueue[3] = 8'b00000000; $display(";A 6685");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6685
            P2_P2_P2_InstQueue[4] = 8'b00000000; $display(";A 6686");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6686
            P2_P2_P2_InstQueue[5] = 8'b00000000; $display(";A 6687");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6687
            P2_P2_P2_InstQueue[6] = 8'b00000000; $display(";A 6688");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6688
            P2_P2_P2_InstQueue[7] = 8'b00000000; $display(";A 6689");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6689
            P2_P2_P2_InstQueue[8] = 8'b00000000; $display(";A 6690");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6690
            P2_P2_P2_InstQueue[9] = 8'b00000000; $display(";A 6691");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6691
            P2_P2_P2_InstQueue[10] = 8'b00000000; $display(";A 6692");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6692
            P2_P2_P2_InstQueue[11] = 8'b00000000; $display(";A 6693");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6693
            P2_P2_P2_InstQueue[12] = 8'b00000000; $display(";A 6694");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6694
            P2_P2_P2_InstQueue[13] = 8'b00000000; $display(";A 6695");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6695
            P2_P2_P2_InstQueue[14] = 8'b00000000; $display(";A 6696");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6696
            P2_P2_P2_InstQueue[15] = 8'b00000000; $display(";A 6697");		//(= P2_P2_P2_InstQueue    0b00000000)) ;6697
            P2_P2_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 6698");		//(= P2_P2_P2_InstQueueRd_Addr    0b00000)) ;6698
            P2_P2_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 6699");		//(= P2_P2_P2_InstQueueWr_Addr    0b00000)) ;6699
            P2_P2_P2_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 6700");		//(= P2_P2_P2_InstAddrPointer    0b00000000000000000000000000000000)) ;6700
            P2_P2_P2_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 6701");		//(= P2_P2_P2_PhyAddrPointer    0b00000000000000000000000000000000)) ;6701
            P2_P2_P2_Extended = 1'b0; $display(";A 6702");		//(= P2_P2_P2_Extended    0b0)) ;6702
            P2_P2_P2_More = 1'b0; $display(";A 6703");		//(= P2_P2_P2_More    0b0)) ;6703
            P2_P2_P2_Flush = 1'b0; $display(";A 6704");		//(= P2_P2_P2_Flush    0b0)) ;6704
            P2_P2_P2_lWord = 16'sb0000000000000000; $display(";A 6705");		//(= P2_P2_P2_lWord    0b0000000000000000)) ;6705
            P2_P2_P2_uWord = 15'sb000000000000000; $display(";A 6706");		//(= P2_P2_P2_uWord    0b000000000000000)) ;6706
            P2_P2_P2_fWord = 32'sb00000000000000000000000000000000; $display(";A 6707");		//(= P2_P2_P2_fWord    0b00000000000000000000000000000000)) ;6707
            P2_P2_P2_CodeFetch <= #1 1'b0; $display(";A 6708");		//(= P2_P2_P2_CodeFetch    0b0)) ;6708
            P2_P2_P2_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 6709");		//(= P2_P2_P2_Datao    0b00000000000000000000000000000000)) ;6709
            P2_P2_P2_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 6710");		//(= P2_P2_P2_EAX    0b00000000000000000000000000000000)) ;6710
            P2_P2_P2_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 6711");		//(= P2_P2_P2_EBX    0b00000000000000000000000000000000)) ;6711
            P2_P2_P2_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 6712");		//(= P2_P2_P2_rEIP    0b00000000000000000000000000000000)) ;6712
            P2_P2_P2_ReadRequest <= #1 1'b0; $display(";A 6713");		//(= P2_P2_P2_ReadRequest    0b0)) ;6713
            P2_P2_P2_MemoryFetch <= #1 1'b0; $display(";A 6714");		//(= P2_P2_P2_MemoryFetch    0b0)) ;6714
            P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6715");		//(= P2_P2_P2_RequestPending    0b0)) ;6715
        end
        else begin
            $display(";A 6680");		//(= (bv-comp P2_P2_P2_RESET  0b1)   0b0)) ;6680
            case (P2_P2_P2_State2)
                4'b0000 :
                    begin
                        $display(";A 6716");		//(= P2_P2_P2_State2    0b0000)) ;6716
                        P2_P2_P2_PhyAddrPointer = P2_P2_P2_rEIP; $display(";A 6717");		//(= P2_P2_P2_PhyAddrPointer    P2_P2_P2_rEIP )) ;6717
                        P2_P2_P2_InstAddrPointer = P2_P2_P2_PhyAddrPointer; $display(";A 6718");		//(= P2_P2_P2_InstAddrPointer    P2_P2_P2_PhyAddrPointer )) ;6718
                        P2_P2_P2_State2 = 4'sb0001; $display(";A 6719");		//(= P2_P2_P2_State2    0b0001)) ;6719
                        P2_P2_P2_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 6720");		//(= P2_P2_P2_rEIP    0b00000000000011111111111111110000)) ;6720
                        P2_P2_P2_ReadRequest <= #1 1'b1; $display(";A 6721");		//(= P2_P2_P2_ReadRequest    0b1)) ;6721
                        P2_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 6722");		//(= P2_P2_P2_MemoryFetch    0b1)) ;6722
                        P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6723");		//(= P2_P2_P2_RequestPending    0b1)) ;6723
                    end
                4'b0001 :
                    begin
                        $display(";A 6724");		//(= P2_P2_P2_State2    0b0001)) ;6724
                        P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6725");		//(= P2_P2_P2_RequestPending    0b1)) ;6725
                        P2_P2_P2_ReadRequest <= #1 1'b1; $display(";A 6726");		//(= P2_P2_P2_ReadRequest    0b1)) ;6726
                        P2_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 6727");		//(= P2_P2_P2_MemoryFetch    0b1)) ;6727
                        P2_P2_P2_CodeFetch <= #1 1'b1; $display(";A 6728");		//(= P2_P2_P2_CodeFetch    0b1)) ;6728
                        if ((P2_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 6729");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6729
                            P2_P2_P2_State2 = 4'sb0010; $display(";A 6731");		//(= P2_P2_P2_State2    0b0010)) ;6731
                        end
                        else begin
                            $display(";A 6730");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6730
                            P2_P2_P2_State2 = 4'sb0001; $display(";A 6732");		//(= P2_P2_P2_State2    0b0001)) ;6732
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 6733");		//(= P2_P2_P2_State2    0b0010)) ;6733
                        P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6734");		//(= P2_P2_P2_RequestPending    0b0)) ;6734
                        P2_P2_P2_InstQueue[P2_P2_P2_InstQueueWr_Addr] = (P2_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 6735");		//(= P2_P2_P2_InstQueue    (bv-smod P2_P2_P2_Datai  0b00000000000000000000000100000000))) ;6735
                        P2_P2_P2_InstQueueWr_Addr = ((P2_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6736");		//(= P2_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6736
                        P2_P2_P2_InstQueue[P2_P2_P2_InstQueueWr_Addr] = (P2_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 6737");		//(= P2_P2_P2_InstQueue    (bv-smod P2_P2_P2_Datai  0b00000000000000000000000100000000))) ;6737
                        P2_P2_P2_InstQueueWr_Addr = ((P2_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6738");		//(= P2_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6738
                        if ((P2_P2_P2_StateBS16 == 1'b1)) begin
                            $display(";A 6739");		//(= (bv-comp P2_P2_P2_StateBS16  0b1)   0b1)) ;6739
                            P2_P2_P2_InstQueue[P2_P2_P2_InstQueueWr_Addr] = ((P2_P2_P2_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 6741");		//(= P2_P2_P2_InstQueue    (bv-smod (bv-sdiv P2_P2_P2_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;6741
                            P2_P2_P2_InstQueueWr_Addr = ((P2_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6742");		//(= P2_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6742
                            P2_P2_P2_InstQueue[P2_P2_P2_InstQueueWr_Addr] = ((P2_P2_P2_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 6743");		//(= P2_P2_P2_InstQueue    (bv-smod (bv-sdiv P2_P2_P2_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;6743
                            P2_P2_P2_InstQueueWr_Addr = ((P2_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6744");		//(= P2_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6744
                            P2_P2_P2_PhyAddrPointer = (P2_P2_P2_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 6745");		//(= P2_P2_P2_PhyAddrPointer    (bv-add P2_P2_P2_PhyAddrPointer  0b00000000000000000000000000000100))) ;6745
                            P2_P2_P2_State2 = 4'sb0101; $display(";A 6746");		//(= P2_P2_P2_State2    0b0101)) ;6746
                        end
                        else begin
                            $display(";A 6740");		//(= (bv-comp P2_P2_P2_StateBS16  0b1)   0b0)) ;6740
                            P2_P2_P2_PhyAddrPointer = (P2_P2_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6747");		//(= P2_P2_P2_PhyAddrPointer    (bv-add P2_P2_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;6747
                            if ((P2_P2_P2_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 6748");		//(= (bool-to-bv (bv-slt P2_P2_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;6748
                                P2_P2_P2_rEIP <= #1 (-P2_P2_P2_PhyAddrPointer); $display(";A 6750");		//(= P2_P2_P2_rEIP    (bv-neg P2_P2_P2_PhyAddrPointer ))) ;6750
                            end
                            else begin
                                $display(";A 6749");		//(= (bool-to-bv (bv-slt P2_P2_P2_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;6749
                                P2_P2_P2_rEIP <= #1 P2_P2_P2_PhyAddrPointer; $display(";A 6751");		//(= P2_P2_P2_rEIP    P2_P2_P2_PhyAddrPointer )) ;6751
                            end
                            P2_P2_P2_State2 = 4'sb0011; $display(";A 6752");		//(= P2_P2_P2_State2    0b0011)) ;6752
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 6753");		//(= P2_P2_P2_State2    0b0011)) ;6753
                        P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6754");		//(= P2_P2_P2_RequestPending    0b1)) ;6754
                        if ((P2_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 6755");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6755
                            P2_P2_P2_State2 = 4'sb0100; $display(";A 6757");		//(= P2_P2_P2_State2    0b0100)) ;6757
                        end
                        else begin
                            $display(";A 6756");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6756
                            P2_P2_P2_State2 = 4'sb0011; $display(";A 6758");		//(= P2_P2_P2_State2    0b0011)) ;6758
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 6759");		//(= P2_P2_P2_State2    0b0100)) ;6759
                        P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6760");		//(= P2_P2_P2_RequestPending    0b0)) ;6760
                        P2_P2_P2_InstQueue[P2_P2_P2_InstQueueWr_Addr] = (P2_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 6761");		//(= P2_P2_P2_InstQueue    (bv-smod P2_P2_P2_Datai  0b00000000000000000000000100000000))) ;6761
                        P2_P2_P2_InstQueueWr_Addr = ((P2_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6762");		//(= P2_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6762
                        P2_P2_P2_InstQueue[P2_P2_P2_InstQueueWr_Addr] = (P2_P2_P2_Datai % 32'b00000000000000000000000100000000); $display(";A 6763");		//(= P2_P2_P2_InstQueue    (bv-smod P2_P2_P2_Datai  0b00000000000000000000000100000000))) ;6763
                        P2_P2_P2_InstQueueWr_Addr = ((P2_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6764");		//(= P2_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6764
                        P2_P2_P2_PhyAddrPointer = (P2_P2_P2_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6765");		//(= P2_P2_P2_PhyAddrPointer    (bv-add P2_P2_P2_PhyAddrPointer  0b00000000000000000000000000000010))) ;6765
                        P2_P2_P2_State2 = 4'sb0101; $display(";A 6766");		//(= P2_P2_P2_State2    0b0101)) ;6766
                    end
                4'b0101 :
                    begin
                        $display(";A 6767");		//(= P2_P2_P2_State2    0b0101)) ;6767
                        case (P2_P2_P2_InstQueue[P2_P2_P2_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 6768");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b10010000)) ;6768
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6769");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6769
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6770");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6770
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6771");		//(= P2_P2_P2_Flush    0b0)) ;6771
                                    P2_P2_P2_More = 1'b0; $display(";A 6772");		//(= P2_P2_P2_More    0b0)) ;6772
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 6773");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b01100110)) ;6773
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6774");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6774
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6775");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6775
                                    P2_P2_P2_Extended = 1'b1; $display(";A 6776");		//(= P2_P2_P2_Extended    0b1)) ;6776
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6777");		//(= P2_P2_P2_Flush    0b0)) ;6777
                                    P2_P2_P2_More = 1'b0; $display(";A 6778");		//(= P2_P2_P2_More    0b0)) ;6778
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 6779");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b11101011)) ;6779
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 6780");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;6780
                                        if ((P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 6782");		//(= (bool-to-bv (bv-gt P2_P2_P2_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;6782
                                            P2_P2_P2_PhyAddrPointer = ((P2_P2_P2_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 6784");		//(= P2_P2_P2_PhyAddrPointer    (bv-sub (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P2_P2_P2_InstQueue 0 )))) ;6784
                                            P2_P2_P2_InstAddrPointer = P2_P2_P2_PhyAddrPointer; $display(";A 6785");		//(= P2_P2_P2_InstAddrPointer    P2_P2_P2_PhyAddrPointer )) ;6785
                                        end
                                        else begin
                                            $display(";A 6783");		//(= (bool-to-bv (bv-gt P2_P2_P2_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;6783
                                            P2_P2_P2_PhyAddrPointer = ((P2_P2_P2_InstAddrPointer + 32'b00000000000000000000000000000010) + P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 6786");		//(= P2_P2_P2_PhyAddrPointer    (bv-add (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000010) P2_P2_P2_InstQueue 0 ))) ;6786
                                            P2_P2_P2_InstAddrPointer = P2_P2_P2_PhyAddrPointer; $display(";A 6787");		//(= P2_P2_P2_InstAddrPointer    P2_P2_P2_PhyAddrPointer )) ;6787
                                        end
                                        P2_P2_P2_Flush = 1'b1; $display(";A 6788");		//(= P2_P2_P2_Flush    0b1)) ;6788
                                        P2_P2_P2_More = 1'b0; $display(";A 6789");		//(= P2_P2_P2_More    0b0)) ;6789
                                    end
                                    else begin
                                        $display(";A 6781");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;6781
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6790");		//(= P2_P2_P2_Flush    0b0)) ;6790
                                        P2_P2_P2_More = 1'b1; $display(";A 6791");		//(= P2_P2_P2_More    0b1)) ;6791
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 6792");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b11101001)) ;6792
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 6793");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;6793
                                        P2_P2_P2_PhyAddrPointer = ((P2_P2_P2_InstAddrPointer + 32'b00000000000000000000000000000101) + P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 6795");		//(= P2_P2_P2_PhyAddrPointer    (bv-add (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000101) P2_P2_P2_InstQueue 0 ))) ;6795
                                        P2_P2_P2_InstAddrPointer = P2_P2_P2_PhyAddrPointer; $display(";A 6796");		//(= P2_P2_P2_InstAddrPointer    P2_P2_P2_PhyAddrPointer )) ;6796
                                        P2_P2_P2_Flush = 1'b1; $display(";A 6797");		//(= P2_P2_P2_Flush    0b1)) ;6797
                                        P2_P2_P2_More = 1'b0; $display(";A 6798");		//(= P2_P2_P2_More    0b0)) ;6798
                                    end
                                    else begin
                                        $display(";A 6794");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;6794
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6799");		//(= P2_P2_P2_Flush    0b0)) ;6799
                                        P2_P2_P2_More = 1'b1; $display(";A 6800");		//(= P2_P2_P2_More    0b1)) ;6800
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 6801");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b11101010)) ;6801
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6802");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6802
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6803");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6803
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6804");		//(= P2_P2_P2_Flush    0b0)) ;6804
                                    P2_P2_P2_More = 1'b0; $display(";A 6805");		//(= P2_P2_P2_More    0b0)) ;6805
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 6806");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b10110000)) ;6806
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6807");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6807
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6808");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6808
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6809");		//(= P2_P2_P2_Flush    0b0)) ;6809
                                    P2_P2_P2_More = 1'b0; $display(";A 6810");		//(= P2_P2_P2_More    0b0)) ;6810
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 6811");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b10111000)) ;6811
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 6812");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;6812
                                        P2_P2_P2_EAX <= #1 ((((P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 6814");		//(= P2_P2_P2_EAX    (bv-add (bv-add (bv-add (bv-mul P2_P2_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P2_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P2_P2_InstQueue 0  0b00000000000000000000000100000000)) P2_P2_P2_InstQueue 0 ))) ;6814
                                        P2_P2_P2_More = 1'b0; $display(";A 6815");		//(= P2_P2_P2_More    0b0)) ;6815
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6816");		//(= P2_P2_P2_Flush    0b0)) ;6816
                                        P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 6817");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;6817
                                        P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 6818");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;6818
                                    end
                                    else begin
                                        $display(";A 6813");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;6813
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6819");		//(= P2_P2_P2_Flush    0b0)) ;6819
                                        P2_P2_P2_More = 1'b1; $display(";A 6820");		//(= P2_P2_P2_More    0b1)) ;6820
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 6821");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b10111011)) ;6821
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 6822");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;6822
                                        P2_P2_P2_EBX <= #1 ((((P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P2_P2_InstQueue[((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 6824");		//(= P2_P2_P2_EBX    (bv-add (bv-add (bv-add (bv-mul P2_P2_P2_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P2_P2_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P2_P2_InstQueue 0  0b00000000000000000000000100000000)) P2_P2_P2_InstQueue 0 ))) ;6824
                                        P2_P2_P2_More = 1'b0; $display(";A 6825");		//(= P2_P2_P2_More    0b0)) ;6825
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6826");		//(= P2_P2_P2_Flush    0b0)) ;6826
                                        P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 6827");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000101))) ;6827
                                        P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 6828");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;6828
                                    end
                                    else begin
                                        $display(";A 6823");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;6823
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6829");		//(= P2_P2_P2_Flush    0b0)) ;6829
                                        P2_P2_P2_More = 1'b1; $display(";A 6830");		//(= P2_P2_P2_More    0b1)) ;6830
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 6831");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b10001011)) ;6831
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6832");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6832
                                        if ((P2_P2_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 6834");		//(= (bool-to-bv (bv-slt P2_P2_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;6834
                                            P2_P2_P2_rEIP <= #1 (-P2_P2_P2_EBX); $display(";A 6836");		//(= P2_P2_P2_rEIP    (bv-neg P2_P2_P2_EBX ))) ;6836
                                        end
                                        else begin
                                            $display(";A 6835");		//(= (bool-to-bv (bv-slt P2_P2_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;6835
                                            P2_P2_P2_rEIP <= #1 P2_P2_P2_EBX; $display(";A 6837");		//(= P2_P2_P2_rEIP    P2_P2_P2_EBX )) ;6837
                                        end
                                        P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6838");		//(= P2_P2_P2_RequestPending    0b1)) ;6838
                                        P2_P2_P2_ReadRequest <= #1 1'b1; $display(";A 6839");		//(= P2_P2_P2_ReadRequest    0b1)) ;6839
                                        P2_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 6840");		//(= P2_P2_P2_MemoryFetch    0b1)) ;6840
                                        P2_P2_P2_CodeFetch <= #1 1'b0; $display(";A 6841");		//(= P2_P2_P2_CodeFetch    0b0)) ;6841
                                        if ((P2_P2_P2_READY_n == 1'b0)) begin
                                            $display(";A 6842");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6842
                                            P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6844");		//(= P2_P2_P2_RequestPending    0b0)) ;6844
                                            P2_P2_P2_uWord = (P2_P2_P2_Datai % 32'b00000000000000001000000000000000); $display(";A 6845");		//(= P2_P2_P2_uWord    (bv-smod P2_P2_P2_Datai  0b00000000000000001000000000000000))) ;6845
                                            if ((P2_P2_P2_StateBS16 == 1'b1)) begin
                                                $display(";A 6846");		//(= (bv-comp P2_P2_P2_StateBS16  0b1)   0b1)) ;6846
                                                P2_P2_P2_lWord = (P2_P2_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 6848");		//(= P2_P2_P2_lWord    (bv-smod P2_P2_P2_Datai  0b00000000000000010000000000000000))) ;6848
                                            end
                                            else begin
                                                $display(";A 6847");		//(= (bv-comp P2_P2_P2_StateBS16  0b1)   0b0)) ;6847
                                                P2_P2_P2_rEIP <= #1 (P2_P2_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 6849");		//(= P2_P2_P2_rEIP    (bv-add P2_P2_P2_rEIP  0b00000000000000000000000000000010))) ;6849
                                                P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6850");		//(= P2_P2_P2_RequestPending    0b1)) ;6850
                                                if ((P2_P2_P2_READY_n == 1'b0)) begin
                                                    $display(";A 6851");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6851
                                                    P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6853");		//(= P2_P2_P2_RequestPending    0b0)) ;6853
                                                    P2_P2_P2_lWord = (P2_P2_P2_Datai % 32'b00000000000000010000000000000000); $display(";A 6854");		//(= P2_P2_P2_lWord    (bv-smod P2_P2_P2_Datai  0b00000000000000010000000000000000))) ;6854
                                                end
                                                else begin
                                                    $display(";A 6852");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6852
                                                end
                                            end
                                            if ((P2_P2_P2_READY_n == 1'b0)) begin
                                                $display(";A 6855");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6855
                                                P2_P2_P2_EAX <= #1 ((P2_P2_P2_uWord * 32'b00000000000000010000000000000000) + P2_P2_P2_lWord); $display(";A 6857");		//(= P2_P2_P2_EAX    (bv-add (bv-mul P2_P2_P2_uWord  0b00000000000000010000000000000000) P2_P2_P2_lWord ))) ;6857
                                                P2_P2_P2_More = 1'b0; $display(";A 6858");		//(= P2_P2_P2_More    0b0)) ;6858
                                                P2_P2_P2_Flush = 1'b0; $display(";A 6859");		//(= P2_P2_P2_Flush    0b0)) ;6859
                                                P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6860");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;6860
                                                P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6861");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6861
                                            end
                                            else begin
                                                $display(";A 6856");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6856
                                            end
                                        end
                                        else begin
                                            $display(";A 6843");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6843
                                        end
                                    end
                                    else begin
                                        $display(";A 6833");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6833
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6862");		//(= P2_P2_P2_Flush    0b0)) ;6862
                                        P2_P2_P2_More = 1'b1; $display(";A 6863");		//(= P2_P2_P2_More    0b1)) ;6863
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 6864");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b10001001)) ;6864
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6865");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6865
                                        if ((P2_P2_P2_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 6867");		//(= (bool-to-bv (bv-slt P2_P2_P2_EBX  0b00000000000000000000000000000000))   0b1)) ;6867
                                            P2_P2_P2_rEIP <= #1 P2_P2_P2_EBX; $display(";A 6869");		//(= P2_P2_P2_rEIP    P2_P2_P2_EBX )) ;6869
                                        end
                                        else begin
                                            $display(";A 6868");		//(= (bool-to-bv (bv-slt P2_P2_P2_EBX  0b00000000000000000000000000000000))   0b0)) ;6868
                                            P2_P2_P2_rEIP <= #1 P2_P2_P2_EBX; $display(";A 6870");		//(= P2_P2_P2_rEIP    P2_P2_P2_EBX )) ;6870
                                        end
                                        P2_P2_P2_lWord = (P2_P2_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 6871");		//(= P2_P2_P2_lWord    (bv-smod P2_P2_P2_EAX  0b00000000000000010000000000000000))) ;6871
                                        P2_P2_P2_uWord = ((P2_P2_P2_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 6872");		//(= P2_P2_P2_uWord    (bv-smod (bv-sdiv P2_P2_P2_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;6872
                                        P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6873");		//(= P2_P2_P2_RequestPending    0b1)) ;6873
                                        P2_P2_P2_ReadRequest <= #1 1'b0; $display(";A 6874");		//(= P2_P2_P2_ReadRequest    0b0)) ;6874
                                        P2_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 6875");		//(= P2_P2_P2_MemoryFetch    0b1)) ;6875
                                        P2_P2_P2_CodeFetch <= #1 1'b0; $display(";A 6876");		//(= P2_P2_P2_CodeFetch    0b0)) ;6876
                                        if (((P2_P2_P2_State == 32'b00000000000000000000000000000010) | (P2_P2_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 6877");		//(= (bv-or (bv-comp P2_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P2_State  0b00000000000000000000000000000100))   0b1)) ;6877
                                            P2_P2_P2_Datao <= #1 ((P2_P2_P2_uWord * 32'b00000000000000010000000000000000) + P2_P2_P2_lWord); $display(";A 6879");		//(= P2_P2_P2_Datao    (bv-add (bv-mul P2_P2_P2_uWord  0b00000000000000010000000000000000) P2_P2_P2_lWord ))) ;6879
                                            if ((P2_P2_P2_READY_n == 1'b0)) begin
                                                $display(";A 6880");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6880
                                                P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6882");		//(= P2_P2_P2_RequestPending    0b0)) ;6882
                                                if ((P2_P2_P2_StateBS16 == 1'b0)) begin
                                                    $display(";A 6883");		//(= (bv-comp P2_P2_P2_StateBS16  0b0)   0b1)) ;6883
                                                    P2_P2_P2_rEIP <= #1 (P2_P2_P2_rEIP + 32'sb00000000000000000000000000000010); $display(";A 6885");		//(= P2_P2_P2_rEIP    (bv-add P2_P2_P2_rEIP  0b00000000000000000000000000000010))) ;6885
                                                    P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6886");		//(= P2_P2_P2_RequestPending    0b1)) ;6886
                                                    P2_P2_P2_ReadRequest <= #1 1'b0; $display(";A 6887");		//(= P2_P2_P2_ReadRequest    0b0)) ;6887
                                                    P2_P2_P2_MemoryFetch <= #1 1'b1; $display(";A 6888");		//(= P2_P2_P2_MemoryFetch    0b1)) ;6888
                                                    P2_P2_P2_CodeFetch <= #1 1'b0; $display(";A 6889");		//(= P2_P2_P2_CodeFetch    0b0)) ;6889
                                                    P2_P2_P2_State2 = 4'sb0110; $display(";A 6890");		//(= P2_P2_P2_State2    0b0110)) ;6890
                                                end
                                                else begin
                                                    $display(";A 6884");		//(= (bv-comp P2_P2_P2_StateBS16  0b0)   0b0)) ;6884
                                                end
                                                P2_P2_P2_More = 1'b0; $display(";A 6891");		//(= P2_P2_P2_More    0b0)) ;6891
                                                P2_P2_P2_Flush = 1'b0; $display(";A 6892");		//(= P2_P2_P2_Flush    0b0)) ;6892
                                                P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6893");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;6893
                                                P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6894");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6894
                                            end
                                            else begin
                                                $display(";A 6881");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6881
                                            end
                                        end
                                        else begin
                                            $display(";A 6878");		//(= (bv-or (bv-comp P2_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P2_State  0b00000000000000000000000000000100))   0b0)) ;6878
                                        end
                                    end
                                    else begin
                                        $display(";A 6866");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6866
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6895");		//(= P2_P2_P2_Flush    0b0)) ;6895
                                        P2_P2_P2_More = 1'b1; $display(";A 6896");		//(= P2_P2_P2_More    0b1)) ;6896
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 6897");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b11100100)) ;6897
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6898");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6898
                                        P2_P2_P2_rEIP <= #1 (P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 6900");		//(= P2_P2_P2_rEIP    (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;6900
                                        P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6901");		//(= P2_P2_P2_RequestPending    0b1)) ;6901
                                        P2_P2_P2_ReadRequest <= #1 1'b1; $display(";A 6902");		//(= P2_P2_P2_ReadRequest    0b1)) ;6902
                                        P2_P2_P2_MemoryFetch <= #1 1'b0; $display(";A 6903");		//(= P2_P2_P2_MemoryFetch    0b0)) ;6903
                                        P2_P2_P2_CodeFetch <= #1 1'b0; $display(";A 6904");		//(= P2_P2_P2_CodeFetch    0b0)) ;6904
                                        if ((P2_P2_P2_READY_n == 1'b0)) begin
                                            $display(";A 6905");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6905
                                            P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6907");		//(= P2_P2_P2_RequestPending    0b0)) ;6907
                                            P2_P2_P2_EAX <= #1 P2_P2_P2_Datai; $display(";A 6908");		//(= P2_P2_P2_EAX    P2_P2_P2_Datai )) ;6908
                                            P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6909");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;6909
                                            P2_P2_P2_InstQueueRd_Addr = (P2_P2_P2_InstQueueRd_Addr + 5'b00010); $display(";A 6910");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-add P2_P2_P2_InstQueueRd_Addr  0b00010))) ;6910
                                            P2_P2_P2_Flush = 1'b0; $display(";A 6911");		//(= P2_P2_P2_Flush    0b0)) ;6911
                                            P2_P2_P2_More = 1'b0; $display(";A 6912");		//(= P2_P2_P2_More    0b0)) ;6912
                                        end
                                        else begin
                                            $display(";A 6906");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6906
                                        end
                                    end
                                    else begin
                                        $display(";A 6899");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6899
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6913");		//(= P2_P2_P2_Flush    0b0)) ;6913
                                        P2_P2_P2_More = 1'b1; $display(";A 6914");		//(= P2_P2_P2_More    0b1)) ;6914
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 6915");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b11100110)) ;6915
                                    if (((P2_P2_P2_InstQueueWr_Addr - P2_P2_P2_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 6916");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;6916
                                        P2_P2_P2_rEIP <= #1 (P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 6918");		//(= P2_P2_P2_rEIP    (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;6918
                                        P2_P2_P2_RequestPending <= #1 1'b1; $display(";A 6919");		//(= P2_P2_P2_RequestPending    0b1)) ;6919
                                        P2_P2_P2_ReadRequest <= #1 1'b0; $display(";A 6920");		//(= P2_P2_P2_ReadRequest    0b0)) ;6920
                                        P2_P2_P2_MemoryFetch <= #1 1'b0; $display(";A 6921");		//(= P2_P2_P2_MemoryFetch    0b0)) ;6921
                                        P2_P2_P2_CodeFetch <= #1 1'b0; $display(";A 6922");		//(= P2_P2_P2_CodeFetch    0b0)) ;6922
                                        if (((P2_P2_P2_State == 32'b00000000000000000000000000000010) | (P2_P2_P2_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 6923");		//(= (bv-or (bv-comp P2_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P2_State  0b00000000000000000000000000000100))   0b1)) ;6923
                                            P2_P2_P2_fWord = (P2_P2_P2_EAX % 32'b00000000000000010000000000000000); $display(";A 6925");		//(= P2_P2_P2_fWord    (bv-smod P2_P2_P2_EAX  0b00000000000000010000000000000000))) ;6925
                                            P2_P2_P2_Datao <= #1 P2_P2_P2_fWord; $display(";A 6926");		//(= P2_P2_P2_Datao    P2_P2_P2_fWord )) ;6926
                                            if ((P2_P2_P2_READY_n == 1'b0)) begin
                                                $display(";A 6927");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6927
                                                P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6929");		//(= P2_P2_P2_RequestPending    0b0)) ;6929
                                                P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6930");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;6930
                                                P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6931");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6931
                                                P2_P2_P2_Flush = 1'b0; $display(";A 6932");		//(= P2_P2_P2_Flush    0b0)) ;6932
                                                P2_P2_P2_More = 1'b0; $display(";A 6933");		//(= P2_P2_P2_More    0b0)) ;6933
                                            end
                                            else begin
                                                $display(";A 6928");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6928
                                            end
                                        end
                                        else begin
                                            $display(";A 6924");		//(= (bv-or (bv-comp P2_P2_P2_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P2_State  0b00000000000000000000000000000100))   0b0)) ;6924
                                        end
                                    end
                                    else begin
                                        $display(";A 6917");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P2_InstQueueWr_Addr  P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;6917
                                        P2_P2_P2_Flush = 1'b0; $display(";A 6934");		//(= P2_P2_P2_Flush    0b0)) ;6934
                                        P2_P2_P2_More = 1'b1; $display(";A 6935");		//(= P2_P2_P2_More    0b1)) ;6935
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 6936");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b00000100)) ;6936
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6937");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6937
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6938");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6938
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6939");		//(= P2_P2_P2_Flush    0b0)) ;6939
                                    P2_P2_P2_More = 1'b0; $display(";A 6940");		//(= P2_P2_P2_More    0b0)) ;6940
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 6941");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b00000101)) ;6941
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6942");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6942
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6943");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6943
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6944");		//(= P2_P2_P2_Flush    0b0)) ;6944
                                    P2_P2_P2_More = 1'b0; $display(";A 6945");		//(= P2_P2_P2_More    0b0)) ;6945
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 6946");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b11010000)) ;6946
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6947");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;6947
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6948");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6948
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6949");		//(= P2_P2_P2_Flush    0b0)) ;6949
                                    P2_P2_P2_More = 1'b0; $display(";A 6950");		//(= P2_P2_P2_More    0b0)) ;6950
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 6951");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b11000000)) ;6951
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 6952");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000010))) ;6952
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 6953");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;6953
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6954");		//(= P2_P2_P2_Flush    0b0)) ;6954
                                    P2_P2_P2_More = 1'b0; $display(";A 6955");		//(= P2_P2_P2_More    0b0)) ;6955
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 6956");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b01000000)) ;6956
                                    P2_P2_P2_EAX <= #1 (P2_P2_P2_EAX + 32'sb00000000000000000000000000000001); $display(";A 6957");		//(= P2_P2_P2_EAX    (bv-add P2_P2_P2_EAX  0b00000000000000000000000000000001))) ;6957
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6958");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6958
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6959");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6959
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6960");		//(= P2_P2_P2_Flush    0b0)) ;6960
                                    P2_P2_P2_More = 1'b0; $display(";A 6961");		//(= P2_P2_P2_More    0b0)) ;6961
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 6962");		//(= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr )   0b01000011)) ;6962
                                    P2_P2_P2_EBX <= #1 (P2_P2_P2_EBX + 32'sb00000000000000000000000000000001); $display(";A 6963");		//(= P2_P2_P2_EBX    (bv-add P2_P2_P2_EBX  0b00000000000000000000000000000001))) ;6963
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6964");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6964
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6965");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6965
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6966");		//(= P2_P2_P2_Flush    0b0)) ;6966
                                    P2_P2_P2_More = 1'b0; $display(";A 6967");		//(= P2_P2_P2_More    0b0)) ;6967
                                end
                            default:
                                begin
                                    $display(";A 6968");		//(= (and (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b10010000) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b01100110) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b11101011) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b11101001) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b11101010) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b10110000) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b10111000) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b10111011) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b10001011) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b10001001) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b11100100) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b11100110) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b00000100) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b00000101) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b11010000) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b11000000) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b01000000) (/= ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ) 0b01000011))   true)) ;6968
                                    P2_P2_P2_InstAddrPointer = (P2_P2_P2_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 6969");		//(= P2_P2_P2_InstAddrPointer    (bv-add P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000001))) ;6969
                                    P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 6970");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;6970
                                    P2_P2_P2_Flush = 1'b0; $display(";A 6971");		//(= P2_P2_P2_Flush    0b0)) ;6971
                                    P2_P2_P2_More = 1'b0; $display(";A 6972");		//(= P2_P2_P2_More    0b0)) ;6972
                                end
                        endcase
                        if (((~(P2_P2_P2_InstQueueRd_Addr < P2_P2_P2_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P2_P2_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P2_P2_P2_Flush) | P2_P2_P2_More))) begin
                            $display(";A 6973");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P2_P2_InstQueueRd_Addr  P2_P2_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P2_P2_Flush ) P2_P2_P2_More ))   0b1)) ;6973
                            P2_P2_P2_State2 = 4'sb0111; $display(";A 6975");		//(= P2_P2_P2_State2    0b0111)) ;6975
                        end
                        else begin
                            $display(";A 6974");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P2_P2_InstQueueRd_Addr  P2_P2_P2_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P2_P2_Flush ) P2_P2_P2_More ))   0b0)) ;6974
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 6976");		//(= P2_P2_P2_State2    0b0110)) ;6976
                        P2_P2_P2_Datao <= #1 ((P2_P2_P2_uWord * 32'b00000000000000010000000000000000) + P2_P2_P2_lWord); $display(";A 6977");		//(= P2_P2_P2_Datao    (bv-add (bv-mul P2_P2_P2_uWord  0b00000000000000010000000000000000) P2_P2_P2_lWord ))) ;6977
                        if ((P2_P2_P2_READY_n == 1'b0)) begin
                            $display(";A 6978");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b1)) ;6978
                            P2_P2_P2_RequestPending <= #1 1'b0; $display(";A 6980");		//(= P2_P2_P2_RequestPending    0b0)) ;6980
                            P2_P2_P2_State2 = 4'sb0101; $display(";A 6981");		//(= P2_P2_P2_State2    0b0101)) ;6981
                        end
                        else begin
                            $display(";A 6979");		//(= (bv-comp P2_P2_P2_READY_n  0b0)   0b0)) ;6979
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 6982");		//(= P2_P2_P2_State2    0b0111)) ;6982
                        if (P2_P2_P2_Flush) begin
                            $display(";A 6983");		//(= P2_P2_P2_Flush    0b1)) ;6983
                            P2_P2_P2_InstQueueRd_Addr = 5'sb00001; $display(";A 6985");		//(= P2_P2_P2_InstQueueRd_Addr    0b00001)) ;6985
                            P2_P2_P2_InstQueueWr_Addr = 5'sb00001; $display(";A 6986");		//(= P2_P2_P2_InstQueueWr_Addr    0b00001)) ;6986
                            if ((P2_P2_P2_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 6987");		//(= (bool-to-bv (bv-slt P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;6987
                                P2_P2_P2_fWord = (-P2_P2_P2_InstAddrPointer); $display(";A 6989");		//(= P2_P2_P2_fWord    (bv-neg P2_P2_P2_InstAddrPointer ))) ;6989
                            end
                            else begin
                                $display(";A 6988");		//(= (bool-to-bv (bv-slt P2_P2_P2_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;6988
                                P2_P2_P2_fWord = P2_P2_P2_InstAddrPointer; $display(";A 6990");		//(= P2_P2_P2_fWord    P2_P2_P2_InstAddrPointer )) ;6990
                            end
                            if (((P2_P2_P2_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 6991");		//(= (bv-comp (bv-smod P2_P2_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;6991
                                P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + (P2_P2_P2_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 6993");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  (bv-smod P2_P2_P2_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;6993
                            end
                            else begin
                                $display(";A 6992");		//(= (bv-comp (bv-smod P2_P2_P2_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;6992
                            end
                        end
                        else begin
                            $display(";A 6984");		//(= P2_P2_P2_Flush    0b0)) ;6984
                        end
                        if (((32'b00000000000000000000000000001111 - P2_P2_P2_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 6994");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;6994
                            P2_P2_P2_State2 = 4'sb1000; $display(";A 6996");		//(= P2_P2_P2_State2    0b1000)) ;6996
                            P2_P2_P2_InstQueueWr_Addr = 5'sb00000; $display(";A 6997");		//(= P2_P2_P2_InstQueueWr_Addr    0b00000)) ;6997
                        end
                        else begin
                            $display(";A 6995");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P2_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;6995
                            P2_P2_P2_State2 = 4'sb1001; $display(";A 6998");		//(= P2_P2_P2_State2    0b1001)) ;6998
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 6999");		//(= P2_P2_P2_State2    0b1000)) ;6999
                        if ((P2_P2_P2_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 7000");		//(= (bool-to-bv (bv-le P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;7000
                            P2_P2_P2_InstQueue[P2_P2_P2_InstQueueWr_Addr] = P2_P2_P2_InstQueue[P2_P2_P2_InstQueueRd_Addr]; $display(";A 7002");		//(= P2_P2_P2_InstQueue    ( P2_P2_P2_InstQueue P2_P2_P2_InstQueueRd_Addr ))) ;7002
                            P2_P2_P2_InstQueueRd_Addr = ((P2_P2_P2_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7003");		//(= P2_P2_P2_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7003
                            P2_P2_P2_InstQueueWr_Addr = ((P2_P2_P2_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7004");		//(= P2_P2_P2_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P2_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7004
                            P2_P2_P2_State2 = 4'sb1000; $display(";A 7005");		//(= P2_P2_P2_State2    0b1000)) ;7005
                        end
                        else begin
                            $display(";A 7001");		//(= (bool-to-bv (bv-le P2_P2_P2_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;7001
                            P2_P2_P2_InstQueueRd_Addr = 5'sb00000; $display(";A 7006");		//(= P2_P2_P2_InstQueueRd_Addr    0b00000)) ;7006
                            P2_P2_P2_State2 = 4'sb1001; $display(";A 7007");		//(= P2_P2_P2_State2    0b1001)) ;7007
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 7008");		//(= P2_P2_P2_State2    0b1001)) ;7008
                        P2_P2_P2_rEIP <= #1 P2_P2_P2_PhyAddrPointer; $display(";A 7009");		//(= P2_P2_P2_rEIP    P2_P2_P2_PhyAddrPointer )) ;7009
                        P2_P2_P2_State2 = 4'sb0001; $display(";A 7010");		//(= P2_P2_P2_State2    0b0001)) ;7010
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:10716
    always @(posedge P2_P2_P2_RESET or posedge P2_P2_P2_CLOCK) begin
        if ((P2_P2_P2_RESET == 1'b1)) begin
            $display(";A 7011");		//(= (bv-comp P2_P2_P2_RESET  0b1)   0b1)) ;7011
            P2_P2_P2_ByteEnable <= #1 4'b0000; $display(";A 7013");		//(= P2_P2_P2_ByteEnable    0b0000)) ;7013
            P2_P2_P2_NonAligned <= #1 1'b0; $display(";A 7014");		//(= P2_P2_P2_NonAligned    0b0)) ;7014
        end
        else begin
            $display(";A 7012");		//(= (bv-comp P2_P2_P2_RESET  0b1)   0b0)) ;7012
            case (P2_P2_P2_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 7015");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000000)) ;7015
                        case ((P2_P2_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 7016");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;7016
                                    P2_P2_P2_ByteEnable <= #1 4'b1110; $display(";A 7017");		//(= P2_P2_P2_ByteEnable    0b1110)) ;7017
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 7018");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;7018
                                    P2_P2_P2_ByteEnable <= #1 4'b1101; $display(";A 7019");		//(= P2_P2_P2_ByteEnable    0b1101)) ;7019
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 7020");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;7020
                                    P2_P2_P2_ByteEnable <= #1 4'b1011; $display(";A 7021");		//(= P2_P2_P2_ByteEnable    0b1011)) ;7021
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 7022");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;7022
                                    P2_P2_P2_ByteEnable <= #1 4'b0111; $display(";A 7023");		//(= P2_P2_P2_ByteEnable    0b0111)) ;7023
                                end
                            default:
                                begin
                                    $display(";A 7024");		//(= (and (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;7024
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 7025");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000001)) ;7025
                        case ((P2_P2_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 7026");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;7026
                                    P2_P2_P2_ByteEnable <= #1 4'b1100; $display(";A 7027");		//(= P2_P2_P2_ByteEnable    0b1100)) ;7027
                                    P2_P2_P2_NonAligned <= #1 1'b0; $display(";A 7028");		//(= P2_P2_P2_NonAligned    0b0)) ;7028
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 7029");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;7029
                                    P2_P2_P2_ByteEnable <= #1 4'b1001; $display(";A 7030");		//(= P2_P2_P2_ByteEnable    0b1001)) ;7030
                                    P2_P2_P2_NonAligned <= #1 1'b0; $display(";A 7031");		//(= P2_P2_P2_NonAligned    0b0)) ;7031
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 7032");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;7032
                                    P2_P2_P2_ByteEnable <= #1 4'b0011; $display(";A 7033");		//(= P2_P2_P2_ByteEnable    0b0011)) ;7033
                                    P2_P2_P2_NonAligned <= #1 1'b0; $display(";A 7034");		//(= P2_P2_P2_NonAligned    0b0)) ;7034
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 7035");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;7035
                                    P2_P2_P2_ByteEnable <= #1 4'b0111; $display(";A 7036");		//(= P2_P2_P2_ByteEnable    0b0111)) ;7036
                                    P2_P2_P2_NonAligned <= #1 1'b1; $display(";A 7037");		//(= P2_P2_P2_NonAligned    0b1)) ;7037
                                end
                            default:
                                begin
                                    $display(";A 7038");		//(= (and (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;7038
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 7039");		//(= P2_P2_P2_DataWidth    0b00000000000000000000000000000010)) ;7039
                        case ((P2_P2_P2_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 7040");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;7040
                                    P2_P2_P2_ByteEnable <= #1 4'b0000; $display(";A 7041");		//(= P2_P2_P2_ByteEnable    0b0000)) ;7041
                                    P2_P2_P2_NonAligned <= #1 1'b0; $display(";A 7042");		//(= P2_P2_P2_NonAligned    0b0)) ;7042
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 7043");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;7043
                                    P2_P2_P2_ByteEnable <= #1 4'b0001; $display(";A 7044");		//(= P2_P2_P2_ByteEnable    0b0001)) ;7044
                                    P2_P2_P2_NonAligned <= #1 1'b1; $display(";A 7045");		//(= P2_P2_P2_NonAligned    0b1)) ;7045
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 7046");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;7046
                                    P2_P2_P2_NonAligned <= #1 1'b1; $display(";A 7047");		//(= P2_P2_P2_NonAligned    0b1)) ;7047
                                    P2_P2_P2_ByteEnable <= #1 4'b0011; $display(";A 7048");		//(= P2_P2_P2_ByteEnable    0b0011)) ;7048
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 7049");		//(= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;7049
                                    P2_P2_P2_NonAligned <= #1 1'b1; $display(";A 7050");		//(= P2_P2_P2_NonAligned    0b1)) ;7050
                                    P2_P2_P2_ByteEnable <= #1 4'b0111; $display(";A 7051");		//(= P2_P2_P2_ByteEnable    0b0111)) ;7051
                                end
                            default:
                                begin
                                    $display(";A 7052");		//(= (and (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P2_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;7052
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 7053");		//(= (and (/= P2_P2_P2_DataWidth  0b00000000000000000000000000000000) (/= P2_P2_P2_DataWidth  0b00000000000000000000000000000001) (/= P2_P2_P2_DataWidth  0b00000000000000000000000000000010))   true)) ;7053
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:10904
    always @(posedge P2_P2_P3_RESET or posedge P2_P2_P3_CLOCK) begin
        if ((P2_P2_P3_RESET == 1'b1)) begin
            $display(";A 7054");		//(= (bv-comp P2_P2_P3_RESET  0b1)   0b1)) ;7054
            P2_P2_P3_BE_n <= #1 4'b0000; $display(";A 7056");		//(= P2_P2_P3_BE_n    0b0000)) ;7056
            P2_P2_P3_Address <= #1 30'sb000000000000000000000000000000; $display(";A 7057");		//(= P2_P2_P3_Address    0b000000000000000000000000000000)) ;7057
            P2_P2_P3_W_R_n <= #1 1'b0; $display(";A 7058");		//(= P2_P2_P3_W_R_n    0b0)) ;7058
            P2_P2_P3_D_C_n <= #1 1'b0; $display(";A 7059");		//(= P2_P2_P3_D_C_n    0b0)) ;7059
            P2_P2_P3_M_IO_n <= #1 1'b0; $display(";A 7060");		//(= P2_P2_P3_M_IO_n    0b0)) ;7060
            P2_P2_P3_ADS_n <= #1 1'b0; $display(";A 7061");		//(= P2_P2_P3_ADS_n    0b0)) ;7061
            P2_P2_P3_State <= #1 3'sb000; $display(";A 7062");		//(= P2_P2_P3_State    0b000)) ;7062
            P2_P2_P3_StateNA <= #1 1'b0; $display(";A 7063");		//(= P2_P2_P3_StateNA    0b0)) ;7063
            P2_P2_P3_StateBS16 <= #1 1'b0; $display(";A 7064");		//(= P2_P2_P3_StateBS16    0b0)) ;7064
            P2_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000000; $display(";A 7065");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000000)) ;7065
        end
        else begin
            $display(";A 7055");		//(= (bv-comp P2_P2_P3_RESET  0b1)   0b0)) ;7055
            case (P2_P2_P3_State)
                3'b000 :
                    begin
                        $display(";A 7066");		//(= P2_P2_P3_State    0b000)) ;7066
                        P2_P2_P3_D_C_n <= #1 1'b1; $display(";A 7067");		//(= P2_P2_P3_D_C_n    0b1)) ;7067
                        P2_P2_P3_ADS_n <= #1 1'b1; $display(";A 7068");		//(= P2_P2_P3_ADS_n    0b1)) ;7068
                        P2_P2_P3_State <= #1 3'sb001; $display(";A 7069");		//(= P2_P2_P3_State    0b001)) ;7069
                        P2_P2_P3_StateNA <= #1 1'b1; $display(";A 7070");		//(= P2_P2_P3_StateNA    0b1)) ;7070
                        P2_P2_P3_StateBS16 <= #1 1'b1; $display(";A 7071");		//(= P2_P2_P3_StateBS16    0b1)) ;7071
                        P2_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 7072");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;7072
                        P2_P2_P3_State <= #1 3'sb001; $display(";A 7073");		//(= P2_P2_P3_State    0b001)) ;7073
                    end
                3'b001 :
                    begin
                        $display(";A 7074");		//(= P2_P2_P3_State    0b001)) ;7074
                        if ((P2_P2_P3_RequestPending == 1'b1)) begin
                            $display(";A 7075");		//(= (bv-comp P2_P2_P3_RequestPending  0b1)   0b1)) ;7075
                            P2_P2_P3_State <= #1 3'sb010; $display(";A 7077");		//(= P2_P2_P3_State    0b010)) ;7077
                        end
                        else begin
                            $display(";A 7076");		//(= (bv-comp P2_P2_P3_RequestPending  0b1)   0b0)) ;7076
                            if ((P2_P2_P3_HOLD == 1'b1)) begin
                                $display(";A 7078");		//(= (bv-comp P2_P2_P3_HOLD  0b1)   0b1)) ;7078
                                P2_P2_P3_State <= #1 3'sb101; $display(";A 7080");		//(= P2_P2_P3_State    0b101)) ;7080
                            end
                            else begin
                                $display(";A 7079");		//(= (bv-comp P2_P2_P3_HOLD  0b1)   0b0)) ;7079
                                P2_P2_P3_State <= #1 3'sb001; $display(";A 7081");		//(= P2_P2_P3_State    0b001)) ;7081
                            end
                        end
                    end
                3'b010 :
                    begin
                        $display(";A 7082");		//(= P2_P2_P3_State    0b010)) ;7082
                        P2_P2_P3_Address <= #1 ((P2_P2_P3_rEIP / 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000000000); $display(";A 7083");		//(= P2_P2_P3_Address    (bv-smod (bv-sdiv P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000))) ;7083
                        P2_P2_P3_BE_n <= #1 P2_P2_P3_ByteEnable; $display(";A 7084");		//(= P2_P2_P3_BE_n    P2_P2_P3_ByteEnable )) ;7084
                        P2_P2_P3_M_IO_n <= #1 P2_P2_P3_MemoryFetch; $display(";A 7085");		//(= P2_P2_P3_M_IO_n    P2_P2_P3_MemoryFetch )) ;7085
                        if ((P2_P2_P3_ReadRequest == 1'b1)) begin
                            $display(";A 7086");		//(= (bv-comp P2_P2_P3_ReadRequest  0b1)   0b1)) ;7086
                            P2_P2_P3_W_R_n <= #1 1'b0; $display(";A 7088");		//(= P2_P2_P3_W_R_n    0b0)) ;7088
                        end
                        else begin
                            $display(";A 7087");		//(= (bv-comp P2_P2_P3_ReadRequest  0b1)   0b0)) ;7087
                            P2_P2_P3_W_R_n <= #1 1'b1; $display(";A 7089");		//(= P2_P2_P3_W_R_n    0b1)) ;7089
                        end
                        if ((P2_P2_P3_CodeFetch == 1'b1)) begin
                            $display(";A 7090");		//(= (bv-comp P2_P2_P3_CodeFetch  0b1)   0b1)) ;7090
                            P2_P2_P3_D_C_n <= #1 1'b0; $display(";A 7092");		//(= P2_P2_P3_D_C_n    0b0)) ;7092
                        end
                        else begin
                            $display(";A 7091");		//(= (bv-comp P2_P2_P3_CodeFetch  0b1)   0b0)) ;7091
                            P2_P2_P3_D_C_n <= #1 1'b1; $display(";A 7093");		//(= P2_P2_P3_D_C_n    0b1)) ;7093
                        end
                        P2_P2_P3_ADS_n <= #1 1'b0; $display(";A 7094");		//(= P2_P2_P3_ADS_n    0b0)) ;7094
                        P2_P2_P3_State <= #1 3'sb011; $display(";A 7095");		//(= P2_P2_P3_State    0b011)) ;7095
                    end
                3'b011 :
                    begin
                        $display(";A 7096");		//(= P2_P2_P3_State    0b011)) ;7096
                        if ((((P2_P2_P3_READY_n == 1'b0) & (P2_P2_P3_HOLD == 1'b0)) & (P2_P2_P3_RequestPending == 1'b1))) begin
                            $display(";A 7097");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b1))   0b1)) ;7097
                            P2_P2_P3_State <= #1 3'sb010; $display(";A 7099");		//(= P2_P2_P3_State    0b010)) ;7099
                        end
                        else begin
                            $display(";A 7098");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b1))   0b0)) ;7098
                            if (((P2_P2_P3_READY_n == 1'b1) & (P2_P2_P3_NA_n == 1'b1))) begin
                                $display(";A 7100");		//(= (bv-and (bv-comp P2_P2_P3_READY_n  0b1) (bv-comp P2_P2_P3_NA_n  0b1))   0b1)) ;7100
                            end
                            else begin
                                $display(";A 7101");		//(= (bv-and (bv-comp P2_P2_P3_READY_n  0b1) (bv-comp P2_P2_P3_NA_n  0b1))   0b0)) ;7101
                                if ((((P2_P2_P3_RequestPending == 1'b1) | (P2_P2_P3_HOLD == 1'b1)) & ((P2_P2_P3_READY_n == 1'b1) & (P2_P2_P3_NA_n == 1'b0)))) begin
                                    $display(";A 7102");		//(= (bv-and (bv-or (bv-comp P2_P2_P3_RequestPending  0b1) (bv-comp P2_P2_P3_HOLD  0b1)) (bv-and (bv-comp P2_P2_P3_READY_n  0b1) (bv-comp P2_P2_P3_NA_n  0b0)))   0b1)) ;7102
                                    P2_P2_P3_State <= #1 3'sb111; $display(";A 7104");		//(= P2_P2_P3_State    0b111)) ;7104
                                end
                                else begin
                                    $display(";A 7103");		//(= (bv-and (bv-or (bv-comp P2_P2_P3_RequestPending  0b1) (bv-comp P2_P2_P3_HOLD  0b1)) (bv-and (bv-comp P2_P2_P3_READY_n  0b1) (bv-comp P2_P2_P3_NA_n  0b0)))   0b0)) ;7103
                                    if (((((P2_P2_P3_RequestPending == 1'b1) & (P2_P2_P3_HOLD == 1'b0)) & (P2_P2_P3_READY_n == 1'b1)) & (P2_P2_P3_NA_n == 1'b0))) begin
                                        $display(";A 7105");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P2_P3_RequestPending  0b1) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_READY_n  0b1)) (bv-comp P2_P2_P3_NA_n  0b0))   0b1)) ;7105
                                        P2_P2_P3_State <= #1 3'sb110; $display(";A 7107");		//(= P2_P2_P3_State    0b110)) ;7107
                                    end
                                    else begin
                                        $display(";A 7106");		//(= (bv-and (bv-and (bv-and (bv-comp P2_P2_P3_RequestPending  0b1) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_READY_n  0b1)) (bv-comp P2_P2_P3_NA_n  0b0))   0b0)) ;7106
                                        if ((((P2_P2_P3_RequestPending == 1'b0) & (P2_P2_P3_HOLD == 1'b0)) & (P2_P2_P3_READY_n == 1'b0))) begin
                                            $display(";A 7108");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_RequestPending  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_READY_n  0b0))   0b1)) ;7108
                                            P2_P2_P3_State <= #1 3'sb001; $display(";A 7110");		//(= P2_P2_P3_State    0b001)) ;7110
                                        end
                                        else begin
                                            $display(";A 7109");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_RequestPending  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_READY_n  0b0))   0b0)) ;7109
                                            if (((P2_P2_P3_HOLD == 1'b1) & (P2_P2_P3_READY_n == 1'b1))) begin
                                                $display(";A 7111");		//(= (bv-and (bv-comp P2_P2_P3_HOLD  0b1) (bv-comp P2_P2_P3_READY_n  0b1))   0b1)) ;7111
                                                P2_P2_P3_State <= #1 3'sb101; $display(";A 7113");		//(= P2_P2_P3_State    0b101)) ;7113
                                            end
                                            else begin
                                                $display(";A 7112");		//(= (bv-and (bv-comp P2_P2_P3_HOLD  0b1) (bv-comp P2_P2_P3_READY_n  0b1))   0b0)) ;7112
                                                P2_P2_P3_State <= #1 3'sb011; $display(";A 7114");		//(= P2_P2_P3_State    0b011)) ;7114
                                            end
                                        end
                                    end
                                end
                            end
                        end
                        P2_P2_P3_StateBS16 <= #1 P2_P2_P3_BS16_n; $display(";A 7115");		//(= P2_P2_P3_StateBS16    P2_P2_P3_BS16_n )) ;7115
                        if ((P2_P2_P3_BS16_n == 1'b0)) begin
                            $display(";A 7116");		//(= (bv-comp P2_P2_P3_BS16_n  0b0)   0b1)) ;7116
                            P2_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 7118");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000001)) ;7118
                        end
                        else begin
                            $display(";A 7117");		//(= (bv-comp P2_P2_P3_BS16_n  0b0)   0b0)) ;7117
                            P2_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 7119");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;7119
                        end
                        P2_P2_P3_StateNA <= #1 P2_P2_P3_NA_n; $display(";A 7120");		//(= P2_P2_P3_StateNA    P2_P2_P3_NA_n )) ;7120
                        P2_P2_P3_ADS_n <= #1 1'b1; $display(";A 7121");		//(= P2_P2_P3_ADS_n    0b1)) ;7121
                    end
                3'b100 :
                    begin
                        $display(";A 7122");		//(= P2_P2_P3_State    0b100)) ;7122
                        if ((((P2_P2_P3_NA_n == 1'b0) & (P2_P2_P3_HOLD == 1'b0)) & (P2_P2_P3_RequestPending == 1'b1))) begin
                            $display(";A 7123");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_NA_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b1))   0b1)) ;7123
                            P2_P2_P3_State <= #1 3'sb110; $display(";A 7125");		//(= P2_P2_P3_State    0b110)) ;7125
                        end
                        else begin
                            $display(";A 7124");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_NA_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b1))   0b0)) ;7124
                            if (((P2_P2_P3_NA_n == 1'b0) & ((P2_P2_P3_HOLD == 1'b1) | (P2_P2_P3_RequestPending == 1'b0)))) begin
                                $display(";A 7126");		//(= (bv-and (bv-comp P2_P2_P3_NA_n  0b0) (bv-or (bv-comp P2_P2_P3_HOLD  0b1) (bv-comp P2_P2_P3_RequestPending  0b0)))   0b1)) ;7126
                                P2_P2_P3_State <= #1 3'sb111; $display(";A 7128");		//(= P2_P2_P3_State    0b111)) ;7128
                            end
                            else begin
                                $display(";A 7127");		//(= (bv-and (bv-comp P2_P2_P3_NA_n  0b0) (bv-or (bv-comp P2_P2_P3_HOLD  0b1) (bv-comp P2_P2_P3_RequestPending  0b0)))   0b0)) ;7127
                                if ((P2_P2_P3_NA_n == 1'b1)) begin
                                    $display(";A 7129");		//(= (bv-comp P2_P2_P3_NA_n  0b1)   0b1)) ;7129
                                    P2_P2_P3_State <= #1 3'sb011; $display(";A 7131");		//(= P2_P2_P3_State    0b011)) ;7131
                                end
                                else begin
                                    $display(";A 7130");		//(= (bv-comp P2_P2_P3_NA_n  0b1)   0b0)) ;7130
                                    P2_P2_P3_State <= #1 3'sb100; $display(";A 7132");		//(= P2_P2_P3_State    0b100)) ;7132
                                end
                            end
                        end
                        P2_P2_P3_StateBS16 <= #1 P2_P2_P3_BS16_n; $display(";A 7133");		//(= P2_P2_P3_StateBS16    P2_P2_P3_BS16_n )) ;7133
                        if ((P2_P2_P3_BS16_n == 1'b0)) begin
                            $display(";A 7134");		//(= (bv-comp P2_P2_P3_BS16_n  0b0)   0b1)) ;7134
                            P2_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000001; $display(";A 7136");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000001)) ;7136
                        end
                        else begin
                            $display(";A 7135");		//(= (bv-comp P2_P2_P3_BS16_n  0b0)   0b0)) ;7135
                            P2_P2_P3_DataWidth <= #1 32'sb00000000000000000000000000000010; $display(";A 7137");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;7137
                        end
                        P2_P2_P3_StateNA <= #1 P2_P2_P3_NA_n; $display(";A 7138");		//(= P2_P2_P3_StateNA    P2_P2_P3_NA_n )) ;7138
                        P2_P2_P3_ADS_n <= #1 1'b1; $display(";A 7139");		//(= P2_P2_P3_ADS_n    0b1)) ;7139
                    end
                3'b101 :
                    begin
                        $display(";A 7140");		//(= P2_P2_P3_State    0b101)) ;7140
                        if (((P2_P2_P3_HOLD == 1'b0) & (P2_P2_P3_RequestPending == 1'b1))) begin
                            $display(";A 7141");		//(= (bv-and (bv-comp P2_P2_P3_HOLD  0b0) (bv-comp P2_P2_P3_RequestPending  0b1))   0b1)) ;7141
                            P2_P2_P3_State <= #1 3'sb010; $display(";A 7143");		//(= P2_P2_P3_State    0b010)) ;7143
                        end
                        else begin
                            $display(";A 7142");		//(= (bv-and (bv-comp P2_P2_P3_HOLD  0b0) (bv-comp P2_P2_P3_RequestPending  0b1))   0b0)) ;7142
                            if (((P2_P2_P3_HOLD == 1'b0) & (P2_P2_P3_RequestPending == 1'b0))) begin
                                $display(";A 7144");		//(= (bv-and (bv-comp P2_P2_P3_HOLD  0b0) (bv-comp P2_P2_P3_RequestPending  0b0))   0b1)) ;7144
                                P2_P2_P3_State <= #1 3'sb001; $display(";A 7146");		//(= P2_P2_P3_State    0b001)) ;7146
                            end
                            else begin
                                $display(";A 7145");		//(= (bv-and (bv-comp P2_P2_P3_HOLD  0b0) (bv-comp P2_P2_P3_RequestPending  0b0))   0b0)) ;7145
                                P2_P2_P3_State <= #1 3'sb101; $display(";A 7147");		//(= P2_P2_P3_State    0b101)) ;7147
                            end
                        end
                    end
                3'b110 :
                    begin
                        $display(";A 7148");		//(= P2_P2_P3_State    0b110)) ;7148
                        P2_P2_P3_Address <= #1 ((P2_P2_P3_rEIP / 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000000000); $display(";A 7149");		//(= P2_P2_P3_Address    (bv-smod (bv-sdiv P2_P2_P3_rEIP  0b00000000000000000000000000000010) 0b00000000000000000000000000000000))) ;7149
                        P2_P2_P3_BE_n <= #1 P2_P2_P3_ByteEnable; $display(";A 7150");		//(= P2_P2_P3_BE_n    P2_P2_P3_ByteEnable )) ;7150
                        P2_P2_P3_M_IO_n <= #1 P2_P2_P3_MemoryFetch; $display(";A 7151");		//(= P2_P2_P3_M_IO_n    P2_P2_P3_MemoryFetch )) ;7151
                        if ((P2_P2_P3_ReadRequest == 1'b1)) begin
                            $display(";A 7152");		//(= (bv-comp P2_P2_P3_ReadRequest  0b1)   0b1)) ;7152
                            P2_P2_P3_W_R_n <= #1 1'b0; $display(";A 7154");		//(= P2_P2_P3_W_R_n    0b0)) ;7154
                        end
                        else begin
                            $display(";A 7153");		//(= (bv-comp P2_P2_P3_ReadRequest  0b1)   0b0)) ;7153
                            P2_P2_P3_W_R_n <= #1 1'b1; $display(";A 7155");		//(= P2_P2_P3_W_R_n    0b1)) ;7155
                        end
                        if ((P2_P2_P3_CodeFetch == 1'b1)) begin
                            $display(";A 7156");		//(= (bv-comp P2_P2_P3_CodeFetch  0b1)   0b1)) ;7156
                            P2_P2_P3_D_C_n <= #1 1'b0; $display(";A 7158");		//(= P2_P2_P3_D_C_n    0b0)) ;7158
                        end
                        else begin
                            $display(";A 7157");		//(= (bv-comp P2_P2_P3_CodeFetch  0b1)   0b0)) ;7157
                            P2_P2_P3_D_C_n <= #1 1'b1; $display(";A 7159");		//(= P2_P2_P3_D_C_n    0b1)) ;7159
                        end
                        P2_P2_P3_ADS_n <= #1 1'b0; $display(";A 7160");		//(= P2_P2_P3_ADS_n    0b0)) ;7160
                        if ((P2_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 7161");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7161
                            P2_P2_P3_State <= #1 3'sb100; $display(";A 7163");		//(= P2_P2_P3_State    0b100)) ;7163
                        end
                        else begin
                            $display(";A 7162");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7162
                            P2_P2_P3_State <= #1 3'sb110; $display(";A 7164");		//(= P2_P2_P3_State    0b110)) ;7164
                        end
                    end
                3'b111 :
                    begin
                        $display(";A 7165");		//(= P2_P2_P3_State    0b111)) ;7165
                        if ((((P2_P2_P3_READY_n == 1'b1) & (P2_P2_P3_RequestPending == 1'b1)) & (P2_P2_P3_HOLD == 1'b0))) begin
                            $display(";A 7166");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b1) (bv-comp P2_P2_P3_RequestPending  0b1)) (bv-comp P2_P2_P3_HOLD  0b0))   0b1)) ;7166
                            P2_P2_P3_State <= #1 3'sb110; $display(";A 7168");		//(= P2_P2_P3_State    0b110)) ;7168
                        end
                        else begin
                            $display(";A 7167");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b1) (bv-comp P2_P2_P3_RequestPending  0b1)) (bv-comp P2_P2_P3_HOLD  0b0))   0b0)) ;7167
                            if (((P2_P2_P3_READY_n == 1'b0) & (P2_P2_P3_HOLD == 1'b1))) begin
                                $display(";A 7169");		//(= (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b1))   0b1)) ;7169
                                P2_P2_P3_State <= #1 3'sb101; $display(";A 7171");		//(= P2_P2_P3_State    0b101)) ;7171
                            end
                            else begin
                                $display(";A 7170");		//(= (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b1))   0b0)) ;7170
                                if ((((P2_P2_P3_READY_n == 1'b0) & (P2_P2_P3_HOLD == 1'b0)) & (P2_P2_P3_RequestPending == 1'b1))) begin
                                    $display(";A 7172");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b1))   0b1)) ;7172
                                    P2_P2_P3_State <= #1 3'sb010; $display(";A 7174");		//(= P2_P2_P3_State    0b010)) ;7174
                                end
                                else begin
                                    $display(";A 7173");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b1))   0b0)) ;7173
                                    if ((((P2_P2_P3_READY_n == 1'b0) & (P2_P2_P3_HOLD == 1'b0)) & (P2_P2_P3_RequestPending == 1'b0))) begin
                                        $display(";A 7175");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b0))   0b1)) ;7175
                                        P2_P2_P3_State <= #1 3'sb001; $display(";A 7177");		//(= P2_P2_P3_State    0b001)) ;7177
                                    end
                                    else begin
                                        $display(";A 7176");		//(= (bv-and (bv-and (bv-comp P2_P2_P3_READY_n  0b0) (bv-comp P2_P2_P3_HOLD  0b0)) (bv-comp P2_P2_P3_RequestPending  0b0))   0b0)) ;7176
                                        P2_P2_P3_State <= #1 3'sb111; $display(";A 7178");		//(= P2_P2_P3_State    0b111)) ;7178
                                    end
                                end
                            end
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:11048
    always @(posedge P2_P2_P3_RESET or posedge P2_P2_P3_CLOCK) begin
        if ((P2_P2_P3_RESET == 1'b1)) begin
            $display(";A 7179");		//(= (bv-comp P2_P2_P3_RESET  0b1)   0b1)) ;7179
            P2_P2_P3_State2 = 4'sb0000; $display(";A 7181");		//(= P2_P2_P3_State2    0b0000)) ;7181
            P2_P2_P3_InstQueue[0] = 8'b00000000; $display(";A 7182");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7182
            P2_P2_P3_InstQueue[1] = 8'b00000000; $display(";A 7183");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7183
            P2_P2_P3_InstQueue[2] = 8'b00000000; $display(";A 7184");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7184
            P2_P2_P3_InstQueue[3] = 8'b00000000; $display(";A 7185");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7185
            P2_P2_P3_InstQueue[4] = 8'b00000000; $display(";A 7186");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7186
            P2_P2_P3_InstQueue[5] = 8'b00000000; $display(";A 7187");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7187
            P2_P2_P3_InstQueue[6] = 8'b00000000; $display(";A 7188");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7188
            P2_P2_P3_InstQueue[7] = 8'b00000000; $display(";A 7189");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7189
            P2_P2_P3_InstQueue[8] = 8'b00000000; $display(";A 7190");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7190
            P2_P2_P3_InstQueue[9] = 8'b00000000; $display(";A 7191");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7191
            P2_P2_P3_InstQueue[10] = 8'b00000000; $display(";A 7192");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7192
            P2_P2_P3_InstQueue[11] = 8'b00000000; $display(";A 7193");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7193
            P2_P2_P3_InstQueue[12] = 8'b00000000; $display(";A 7194");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7194
            P2_P2_P3_InstQueue[13] = 8'b00000000; $display(";A 7195");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7195
            P2_P2_P3_InstQueue[14] = 8'b00000000; $display(";A 7196");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7196
            P2_P2_P3_InstQueue[15] = 8'b00000000; $display(";A 7197");		//(= P2_P2_P3_InstQueue    0b00000000)) ;7197
            P2_P2_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 7198");		//(= P2_P2_P3_InstQueueRd_Addr    0b00000)) ;7198
            P2_P2_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 7199");		//(= P2_P2_P3_InstQueueWr_Addr    0b00000)) ;7199
            P2_P2_P3_InstAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 7200");		//(= P2_P2_P3_InstAddrPointer    0b00000000000000000000000000000000)) ;7200
            P2_P2_P3_PhyAddrPointer = 32'sb00000000000000000000000000000000; $display(";A 7201");		//(= P2_P2_P3_PhyAddrPointer    0b00000000000000000000000000000000)) ;7201
            P2_P2_P3_Extended = 1'b0; $display(";A 7202");		//(= P2_P2_P3_Extended    0b0)) ;7202
            P2_P2_P3_More = 1'b0; $display(";A 7203");		//(= P2_P2_P3_More    0b0)) ;7203
            P2_P2_P3_Flush = 1'b0; $display(";A 7204");		//(= P2_P2_P3_Flush    0b0)) ;7204
            P2_P2_P3_lWord = 16'sb0000000000000000; $display(";A 7205");		//(= P2_P2_P3_lWord    0b0000000000000000)) ;7205
            P2_P2_P3_uWord = 15'sb000000000000000; $display(";A 7206");		//(= P2_P2_P3_uWord    0b000000000000000)) ;7206
            P2_P2_P3_fWord = 32'sb00000000000000000000000000000000; $display(";A 7207");		//(= P2_P2_P3_fWord    0b00000000000000000000000000000000)) ;7207
            P2_P2_P3_CodeFetch <= #1 1'b0; $display(";A 7208");		//(= P2_P2_P3_CodeFetch    0b0)) ;7208
            P2_P2_P3_Datao <= #1 32'sb00000000000000000000000000000000; $display(";A 7209");		//(= P2_P2_P3_Datao    0b00000000000000000000000000000000)) ;7209
            P2_P2_P3_EAX <= #1 32'sb00000000000000000000000000000000; $display(";A 7210");		//(= P2_P2_P3_EAX    0b00000000000000000000000000000000)) ;7210
            P2_P2_P3_EBX <= #1 32'sb00000000000000000000000000000000; $display(";A 7211");		//(= P2_P2_P3_EBX    0b00000000000000000000000000000000)) ;7211
            P2_P2_P3_rEIP <= #1 32'sb00000000000000000000000000000000; $display(";A 7212");		//(= P2_P2_P3_rEIP    0b00000000000000000000000000000000)) ;7212
            P2_P2_P3_ReadRequest <= #1 1'b0; $display(";A 7213");		//(= P2_P2_P3_ReadRequest    0b0)) ;7213
            P2_P2_P3_MemoryFetch <= #1 1'b0; $display(";A 7214");		//(= P2_P2_P3_MemoryFetch    0b0)) ;7214
            P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7215");		//(= P2_P2_P3_RequestPending    0b0)) ;7215
        end
        else begin
            $display(";A 7180");		//(= (bv-comp P2_P2_P3_RESET  0b1)   0b0)) ;7180
            case (P2_P2_P3_State2)
                4'b0000 :
                    begin
                        $display(";A 7216");		//(= P2_P2_P3_State2    0b0000)) ;7216
                        P2_P2_P3_PhyAddrPointer = P2_P2_P3_rEIP; $display(";A 7217");		//(= P2_P2_P3_PhyAddrPointer    P2_P2_P3_rEIP )) ;7217
                        P2_P2_P3_InstAddrPointer = P2_P2_P3_PhyAddrPointer; $display(";A 7218");		//(= P2_P2_P3_InstAddrPointer    P2_P2_P3_PhyAddrPointer )) ;7218
                        P2_P2_P3_State2 = 4'sb0001; $display(";A 7219");		//(= P2_P2_P3_State2    0b0001)) ;7219
                        P2_P2_P3_rEIP <= #1 32'b00000000000011111111111111110000; $display(";A 7220");		//(= P2_P2_P3_rEIP    0b00000000000011111111111111110000)) ;7220
                        P2_P2_P3_ReadRequest <= #1 1'b1; $display(";A 7221");		//(= P2_P2_P3_ReadRequest    0b1)) ;7221
                        P2_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 7222");		//(= P2_P2_P3_MemoryFetch    0b1)) ;7222
                        P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7223");		//(= P2_P2_P3_RequestPending    0b1)) ;7223
                    end
                4'b0001 :
                    begin
                        $display(";A 7224");		//(= P2_P2_P3_State2    0b0001)) ;7224
                        P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7225");		//(= P2_P2_P3_RequestPending    0b1)) ;7225
                        P2_P2_P3_ReadRequest <= #1 1'b1; $display(";A 7226");		//(= P2_P2_P3_ReadRequest    0b1)) ;7226
                        P2_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 7227");		//(= P2_P2_P3_MemoryFetch    0b1)) ;7227
                        P2_P2_P3_CodeFetch <= #1 1'b1; $display(";A 7228");		//(= P2_P2_P3_CodeFetch    0b1)) ;7228
                        if ((P2_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 7229");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7229
                            P2_P2_P3_State2 = 4'sb0010; $display(";A 7231");		//(= P2_P2_P3_State2    0b0010)) ;7231
                        end
                        else begin
                            $display(";A 7230");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7230
                            P2_P2_P3_State2 = 4'sb0001; $display(";A 7232");		//(= P2_P2_P3_State2    0b0001)) ;7232
                        end
                    end
                4'b0010 :
                    begin
                        $display(";A 7233");		//(= P2_P2_P3_State2    0b0010)) ;7233
                        P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7234");		//(= P2_P2_P3_RequestPending    0b0)) ;7234
                        P2_P2_P3_InstQueue[P2_P2_P3_InstQueueWr_Addr] = (P2_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 7235");		//(= P2_P2_P3_InstQueue    (bv-smod P2_P2_P3_Datai  0b00000000000000000000000100000000))) ;7235
                        P2_P2_P3_InstQueueWr_Addr = ((P2_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7236");		//(= P2_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7236
                        P2_P2_P3_InstQueue[P2_P2_P3_InstQueueWr_Addr] = (P2_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 7237");		//(= P2_P2_P3_InstQueue    (bv-smod P2_P2_P3_Datai  0b00000000000000000000000100000000))) ;7237
                        P2_P2_P3_InstQueueWr_Addr = ((P2_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7238");		//(= P2_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7238
                        if ((P2_P2_P3_StateBS16 == 1'b1)) begin
                            $display(";A 7239");		//(= (bv-comp P2_P2_P3_StateBS16  0b1)   0b1)) ;7239
                            P2_P2_P3_InstQueue[P2_P2_P3_InstQueueWr_Addr] = ((P2_P2_P3_Datai / 32'b00000000000000010000000000000000) % 32'b00000000000000000000000100000000); $display(";A 7241");		//(= P2_P2_P3_InstQueue    (bv-smod (bv-sdiv P2_P2_P3_Datai  0b00000000000000010000000000000000) 0b00000000000000000000000100000000))) ;7241
                            P2_P2_P3_InstQueueWr_Addr = ((P2_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7242");		//(= P2_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7242
                            P2_P2_P3_InstQueue[P2_P2_P3_InstQueueWr_Addr] = ((P2_P2_P3_Datai / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000100000000); $display(";A 7243");		//(= P2_P2_P3_InstQueue    (bv-smod (bv-sdiv P2_P2_P3_Datai  0b00000001000000000000000000000000) 0b00000000000000000000000100000000))) ;7243
                            P2_P2_P3_InstQueueWr_Addr = ((P2_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7244");		//(= P2_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7244
                            P2_P2_P3_PhyAddrPointer = (P2_P2_P3_PhyAddrPointer + 32'sb00000000000000000000000000000100); $display(";A 7245");		//(= P2_P2_P3_PhyAddrPointer    (bv-add P2_P2_P3_PhyAddrPointer  0b00000000000000000000000000000100))) ;7245
                            P2_P2_P3_State2 = 4'sb0101; $display(";A 7246");		//(= P2_P2_P3_State2    0b0101)) ;7246
                        end
                        else begin
                            $display(";A 7240");		//(= (bv-comp P2_P2_P3_StateBS16  0b1)   0b0)) ;7240
                            P2_P2_P3_PhyAddrPointer = (P2_P2_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7247");		//(= P2_P2_P3_PhyAddrPointer    (bv-add P2_P2_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;7247
                            if ((P2_P2_P3_PhyAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 7248");		//(= (bool-to-bv (bv-slt P2_P2_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b1)) ;7248
                                P2_P2_P3_rEIP <= #1 (-P2_P2_P3_PhyAddrPointer); $display(";A 7250");		//(= P2_P2_P3_rEIP    (bv-neg P2_P2_P3_PhyAddrPointer ))) ;7250
                            end
                            else begin
                                $display(";A 7249");		//(= (bool-to-bv (bv-slt P2_P2_P3_PhyAddrPointer  0b00000000000000000000000000000000))   0b0)) ;7249
                                P2_P2_P3_rEIP <= #1 P2_P2_P3_PhyAddrPointer; $display(";A 7251");		//(= P2_P2_P3_rEIP    P2_P2_P3_PhyAddrPointer )) ;7251
                            end
                            P2_P2_P3_State2 = 4'sb0011; $display(";A 7252");		//(= P2_P2_P3_State2    0b0011)) ;7252
                        end
                    end
                4'b0011 :
                    begin
                        $display(";A 7253");		//(= P2_P2_P3_State2    0b0011)) ;7253
                        P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7254");		//(= P2_P2_P3_RequestPending    0b1)) ;7254
                        if ((P2_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 7255");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7255
                            P2_P2_P3_State2 = 4'sb0100; $display(";A 7257");		//(= P2_P2_P3_State2    0b0100)) ;7257
                        end
                        else begin
                            $display(";A 7256");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7256
                            P2_P2_P3_State2 = 4'sb0011; $display(";A 7258");		//(= P2_P2_P3_State2    0b0011)) ;7258
                        end
                    end
                4'b0100 :
                    begin
                        $display(";A 7259");		//(= P2_P2_P3_State2    0b0100)) ;7259
                        P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7260");		//(= P2_P2_P3_RequestPending    0b0)) ;7260
                        P2_P2_P3_InstQueue[P2_P2_P3_InstQueueWr_Addr] = (P2_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 7261");		//(= P2_P2_P3_InstQueue    (bv-smod P2_P2_P3_Datai  0b00000000000000000000000100000000))) ;7261
                        P2_P2_P3_InstQueueWr_Addr = ((P2_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7262");		//(= P2_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7262
                        P2_P2_P3_InstQueue[P2_P2_P3_InstQueueWr_Addr] = (P2_P2_P3_Datai % 32'b00000000000000000000000100000000); $display(";A 7263");		//(= P2_P2_P3_InstQueue    (bv-smod P2_P2_P3_Datai  0b00000000000000000000000100000000))) ;7263
                        P2_P2_P3_InstQueueWr_Addr = ((P2_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7264");		//(= P2_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7264
                        P2_P2_P3_PhyAddrPointer = (P2_P2_P3_PhyAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7265");		//(= P2_P2_P3_PhyAddrPointer    (bv-add P2_P2_P3_PhyAddrPointer  0b00000000000000000000000000000010))) ;7265
                        P2_P2_P3_State2 = 4'sb0101; $display(";A 7266");		//(= P2_P2_P3_State2    0b0101)) ;7266
                    end
                4'b0101 :
                    begin
                        $display(";A 7267");		//(= P2_P2_P3_State2    0b0101)) ;7267
                        case (P2_P2_P3_InstQueue[P2_P2_P3_InstQueueRd_Addr])
                            8'b10010000 :
                                begin
                                    $display(";A 7268");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b10010000)) ;7268
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7269");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7269
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7270");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7270
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7271");		//(= P2_P2_P3_Flush    0b0)) ;7271
                                    P2_P2_P3_More = 1'b0; $display(";A 7272");		//(= P2_P2_P3_More    0b0)) ;7272
                                end
                            8'b01100110 :
                                begin
                                    $display(";A 7273");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b01100110)) ;7273
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7274");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7274
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7275");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7275
                                    P2_P2_P3_Extended = 1'b1; $display(";A 7276");		//(= P2_P2_P3_Extended    0b1)) ;7276
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7277");		//(= P2_P2_P3_Flush    0b0)) ;7277
                                    P2_P2_P3_More = 1'b0; $display(";A 7278");		//(= P2_P2_P3_More    0b0)) ;7278
                                end
                            8'b11101011 :
                                begin
                                    $display(";A 7279");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b11101011)) ;7279
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000011)) begin
                                        $display(";A 7280");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;7280
                                        if ((P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)] > 32'b00000000000000000000000001111111)) begin
                                            $display(";A 7282");		//(= (bool-to-bv (bv-gt P2_P2_P3_InstQueue 0  0b00000000000000000000000001111111))   0b1)) ;7282
                                            P2_P2_P3_PhyAddrPointer = ((P2_P2_P3_InstAddrPointer + 32'b00000000000000000000000000000001) - (32'b00000000000000000000000011111111 - P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)])); $display(";A 7284");		//(= P2_P2_P3_PhyAddrPointer    (bv-sub (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001) (bv-sub 0b00000000000000000000000011111111 P2_P2_P3_InstQueue 0 )))) ;7284
                                            P2_P2_P3_InstAddrPointer = P2_P2_P3_PhyAddrPointer; $display(";A 7285");		//(= P2_P2_P3_InstAddrPointer    P2_P2_P3_PhyAddrPointer )) ;7285
                                        end
                                        else begin
                                            $display(";A 7283");		//(= (bool-to-bv (bv-gt P2_P2_P3_InstQueue 0  0b00000000000000000000000001111111))   0b0)) ;7283
                                            P2_P2_P3_PhyAddrPointer = ((P2_P2_P3_InstAddrPointer + 32'b00000000000000000000000000000010) + P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 7286");		//(= P2_P2_P3_PhyAddrPointer    (bv-add (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000010) P2_P2_P3_InstQueue 0 ))) ;7286
                                            P2_P2_P3_InstAddrPointer = P2_P2_P3_PhyAddrPointer; $display(";A 7287");		//(= P2_P2_P3_InstAddrPointer    P2_P2_P3_PhyAddrPointer )) ;7287
                                        end
                                        P2_P2_P3_Flush = 1'b1; $display(";A 7288");		//(= P2_P2_P3_Flush    0b1)) ;7288
                                        P2_P2_P3_More = 1'b0; $display(";A 7289");		//(= P2_P2_P3_More    0b0)) ;7289
                                    end
                                    else begin
                                        $display(";A 7281");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;7281
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7290");		//(= P2_P2_P3_Flush    0b0)) ;7290
                                        P2_P2_P3_More = 1'b1; $display(";A 7291");		//(= P2_P2_P3_More    0b1)) ;7291
                                    end
                                end
                            8'b11101001 :
                                begin
                                    $display(";A 7292");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b11101001)) ;7292
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 7293");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;7293
                                        P2_P2_P3_PhyAddrPointer = ((P2_P2_P3_InstAddrPointer + 32'b00000000000000000000000000000101) + P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 7295");		//(= P2_P2_P3_PhyAddrPointer    (bv-add (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000101) P2_P2_P3_InstQueue 0 ))) ;7295
                                        P2_P2_P3_InstAddrPointer = P2_P2_P3_PhyAddrPointer; $display(";A 7296");		//(= P2_P2_P3_InstAddrPointer    P2_P2_P3_PhyAddrPointer )) ;7296
                                        P2_P2_P3_Flush = 1'b1; $display(";A 7297");		//(= P2_P2_P3_Flush    0b1)) ;7297
                                        P2_P2_P3_More = 1'b0; $display(";A 7298");		//(= P2_P2_P3_More    0b0)) ;7298
                                    end
                                    else begin
                                        $display(";A 7294");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;7294
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7299");		//(= P2_P2_P3_Flush    0b0)) ;7299
                                        P2_P2_P3_More = 1'b1; $display(";A 7300");		//(= P2_P2_P3_More    0b1)) ;7300
                                    end
                                end
                            8'b11101010 :
                                begin
                                    $display(";A 7301");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b11101010)) ;7301
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7302");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7302
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7303");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7303
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7304");		//(= P2_P2_P3_Flush    0b0)) ;7304
                                    P2_P2_P3_More = 1'b0; $display(";A 7305");		//(= P2_P2_P3_More    0b0)) ;7305
                                end
                            8'b10110000 :
                                begin
                                    $display(";A 7306");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b10110000)) ;7306
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7307");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7307
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7308");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7308
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7309");		//(= P2_P2_P3_Flush    0b0)) ;7309
                                    P2_P2_P3_More = 1'b0; $display(";A 7310");		//(= P2_P2_P3_More    0b0)) ;7310
                                end
                            8'b10111000 :
                                begin
                                    $display(";A 7311");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b10111000)) ;7311
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 7312");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;7312
                                        P2_P2_P3_EAX <= #1 ((((P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000)]); $display(";A 7314");		//(= P2_P2_P3_EAX    (bv-add (bv-add (bv-add (bv-mul P2_P2_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P2_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P2_P3_InstQueue 0  0b00000000000000000000000100000000)) P2_P2_P3_InstQueue 0 ))) ;7314
                                        P2_P2_P3_More = 1'b0; $display(";A 7315");		//(= P2_P2_P3_More    0b0)) ;7315
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7316");		//(= P2_P2_P3_Flush    0b0)) ;7316
                                        P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 7317");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;7317
                                        P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 7318");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;7318
                                    end
                                    else begin
                                        $display(";A 7313");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;7313
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7319");		//(= P2_P2_P3_Flush    0b0)) ;7319
                                        P2_P2_P3_More = 1'b1; $display(";A 7320");		//(= P2_P2_P3_More    0b1)) ;7320
                                    end
                                end
                            8'b10111011 :
                                begin
                                    $display(";A 7321");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b10111011)) ;7321
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000101)) begin
                                        $display(";A 7322");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b1)) ;7322
                                        P2_P2_P3_EBX <= #1 ((((P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000100) % 32'b00000000000000000000000000010000)] * 32'b00000000100000000000000000000000) + (P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000011) % 32'b00000000000000000000000000010000)] * 32'b00000000000000010000000000000000)) + (P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000)] * 32'b00000000000000000000000100000000)) + P2_P2_P3_InstQueue[((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000000001)]); $display(";A 7324");		//(= P2_P2_P3_EBX    (bv-add (bv-add (bv-add (bv-mul P2_P2_P3_InstQueue 0  0b00000000100000000000000000000000) (bv-mul P2_P2_P3_InstQueue 0  0b00000000000000010000000000000000)) (bv-mul P2_P2_P3_InstQueue 0  0b00000000000000000000000100000000)) P2_P2_P3_InstQueue 0 ))) ;7324
                                        P2_P2_P3_More = 1'b0; $display(";A 7325");		//(= P2_P2_P3_More    0b0)) ;7325
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7326");		//(= P2_P2_P3_Flush    0b0)) ;7326
                                        P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000101); $display(";A 7327");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000101))) ;7327
                                        P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000101) % 32'b00000000000000000000000000010000); $display(";A 7328");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000101) 0b00000000000000000000000000010000))) ;7328
                                    end
                                    else begin
                                        $display(";A 7323");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000101))   0b0)) ;7323
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7329");		//(= P2_P2_P3_Flush    0b0)) ;7329
                                        P2_P2_P3_More = 1'b1; $display(";A 7330");		//(= P2_P2_P3_More    0b1)) ;7330
                                    end
                                end
                            8'b10001011 :
                                begin
                                    $display(";A 7331");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b10001011)) ;7331
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 7332");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;7332
                                        if ((P2_P2_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 7334");		//(= (bool-to-bv (bv-slt P2_P2_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;7334
                                            P2_P2_P3_rEIP <= #1 (-P2_P2_P3_EBX); $display(";A 7336");		//(= P2_P2_P3_rEIP    (bv-neg P2_P2_P3_EBX ))) ;7336
                                        end
                                        else begin
                                            $display(";A 7335");		//(= (bool-to-bv (bv-slt P2_P2_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;7335
                                            P2_P2_P3_rEIP <= #1 P2_P2_P3_EBX; $display(";A 7337");		//(= P2_P2_P3_rEIP    P2_P2_P3_EBX )) ;7337
                                        end
                                        P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7338");		//(= P2_P2_P3_RequestPending    0b1)) ;7338
                                        P2_P2_P3_ReadRequest <= #1 1'b1; $display(";A 7339");		//(= P2_P2_P3_ReadRequest    0b1)) ;7339
                                        P2_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 7340");		//(= P2_P2_P3_MemoryFetch    0b1)) ;7340
                                        P2_P2_P3_CodeFetch <= #1 1'b0; $display(";A 7341");		//(= P2_P2_P3_CodeFetch    0b0)) ;7341
                                        if ((P2_P2_P3_READY_n == 1'b0)) begin
                                            $display(";A 7342");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7342
                                            P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7344");		//(= P2_P2_P3_RequestPending    0b0)) ;7344
                                            P2_P2_P3_uWord = (P2_P2_P3_Datai % 32'b00000000000000001000000000000000); $display(";A 7345");		//(= P2_P2_P3_uWord    (bv-smod P2_P2_P3_Datai  0b00000000000000001000000000000000))) ;7345
                                            if ((P2_P2_P3_StateBS16 == 1'b1)) begin
                                                $display(";A 7346");		//(= (bv-comp P2_P2_P3_StateBS16  0b1)   0b1)) ;7346
                                                P2_P2_P3_lWord = (P2_P2_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 7348");		//(= P2_P2_P3_lWord    (bv-smod P2_P2_P3_Datai  0b00000000000000010000000000000000))) ;7348
                                            end
                                            else begin
                                                $display(";A 7347");		//(= (bv-comp P2_P2_P3_StateBS16  0b1)   0b0)) ;7347
                                                P2_P2_P3_rEIP <= #1 (P2_P2_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 7349");		//(= P2_P2_P3_rEIP    (bv-add P2_P2_P3_rEIP  0b00000000000000000000000000000010))) ;7349
                                                P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7350");		//(= P2_P2_P3_RequestPending    0b1)) ;7350
                                                if ((P2_P2_P3_READY_n == 1'b0)) begin
                                                    $display(";A 7351");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7351
                                                    P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7353");		//(= P2_P2_P3_RequestPending    0b0)) ;7353
                                                    P2_P2_P3_lWord = (P2_P2_P3_Datai % 32'b00000000000000010000000000000000); $display(";A 7354");		//(= P2_P2_P3_lWord    (bv-smod P2_P2_P3_Datai  0b00000000000000010000000000000000))) ;7354
                                                end
                                                else begin
                                                    $display(";A 7352");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7352
                                                end
                                            end
                                            if ((P2_P2_P3_READY_n == 1'b0)) begin
                                                $display(";A 7355");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7355
                                                P2_P2_P3_EAX <= #1 ((P2_P2_P3_uWord * 32'b00000000000000010000000000000000) + P2_P2_P3_lWord); $display(";A 7357");		//(= P2_P2_P3_EAX    (bv-add (bv-mul P2_P2_P3_uWord  0b00000000000000010000000000000000) P2_P2_P3_lWord ))) ;7357
                                                P2_P2_P3_More = 1'b0; $display(";A 7358");		//(= P2_P2_P3_More    0b0)) ;7358
                                                P2_P2_P3_Flush = 1'b0; $display(";A 7359");		//(= P2_P2_P3_Flush    0b0)) ;7359
                                                P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7360");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;7360
                                                P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 7361");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;7361
                                            end
                                            else begin
                                                $display(";A 7356");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7356
                                            end
                                        end
                                        else begin
                                            $display(";A 7343");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7343
                                        end
                                    end
                                    else begin
                                        $display(";A 7333");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;7333
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7362");		//(= P2_P2_P3_Flush    0b0)) ;7362
                                        P2_P2_P3_More = 1'b1; $display(";A 7363");		//(= P2_P2_P3_More    0b1)) ;7363
                                    end
                                end
                            8'b10001001 :
                                begin
                                    $display(";A 7364");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b10001001)) ;7364
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 7365");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;7365
                                        if ((P2_P2_P3_EBX < 32'sb00000000000000000000000000000000)) begin
                                            $display(";A 7367");		//(= (bool-to-bv (bv-slt P2_P2_P3_EBX  0b00000000000000000000000000000000))   0b1)) ;7367
                                            P2_P2_P3_rEIP <= #1 P2_P2_P3_EBX; $display(";A 7369");		//(= P2_P2_P3_rEIP    P2_P2_P3_EBX )) ;7369
                                        end
                                        else begin
                                            $display(";A 7368");		//(= (bool-to-bv (bv-slt P2_P2_P3_EBX  0b00000000000000000000000000000000))   0b0)) ;7368
                                            P2_P2_P3_rEIP <= #1 P2_P2_P3_EBX; $display(";A 7370");		//(= P2_P2_P3_rEIP    P2_P2_P3_EBX )) ;7370
                                        end
                                        P2_P2_P3_lWord = (P2_P2_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 7371");		//(= P2_P2_P3_lWord    (bv-smod P2_P2_P3_EAX  0b00000000000000010000000000000000))) ;7371
                                        P2_P2_P3_uWord = ((P2_P2_P3_EAX / 32'b00000000000000010000000000000000) % 32'b00000000000000001000000000000000); $display(";A 7372");		//(= P2_P2_P3_uWord    (bv-smod (bv-sdiv P2_P2_P3_EAX  0b00000000000000010000000000000000) 0b00000000000000001000000000000000))) ;7372
                                        P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7373");		//(= P2_P2_P3_RequestPending    0b1)) ;7373
                                        P2_P2_P3_ReadRequest <= #1 1'b0; $display(";A 7374");		//(= P2_P2_P3_ReadRequest    0b0)) ;7374
                                        P2_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 7375");		//(= P2_P2_P3_MemoryFetch    0b1)) ;7375
                                        P2_P2_P3_CodeFetch <= #1 1'b0; $display(";A 7376");		//(= P2_P2_P3_CodeFetch    0b0)) ;7376
                                        if (((P2_P2_P3_State == 32'b00000000000000000000000000000010) | (P2_P2_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 7377");		//(= (bv-or (bv-comp P2_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P3_State  0b00000000000000000000000000000100))   0b1)) ;7377
                                            P2_P2_P3_Datao <= #1 ((P2_P2_P3_uWord * 32'b00000000000000010000000000000000) + P2_P2_P3_lWord); $display(";A 7379");		//(= P2_P2_P3_Datao    (bv-add (bv-mul P2_P2_P3_uWord  0b00000000000000010000000000000000) P2_P2_P3_lWord ))) ;7379
                                            if ((P2_P2_P3_READY_n == 1'b0)) begin
                                                $display(";A 7380");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7380
                                                P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7382");		//(= P2_P2_P3_RequestPending    0b0)) ;7382
                                                if ((P2_P2_P3_StateBS16 == 1'b0)) begin
                                                    $display(";A 7383");		//(= (bv-comp P2_P2_P3_StateBS16  0b0)   0b1)) ;7383
                                                    P2_P2_P3_rEIP <= #1 (P2_P2_P3_rEIP + 32'sb00000000000000000000000000000010); $display(";A 7385");		//(= P2_P2_P3_rEIP    (bv-add P2_P2_P3_rEIP  0b00000000000000000000000000000010))) ;7385
                                                    P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7386");		//(= P2_P2_P3_RequestPending    0b1)) ;7386
                                                    P2_P2_P3_ReadRequest <= #1 1'b0; $display(";A 7387");		//(= P2_P2_P3_ReadRequest    0b0)) ;7387
                                                    P2_P2_P3_MemoryFetch <= #1 1'b1; $display(";A 7388");		//(= P2_P2_P3_MemoryFetch    0b1)) ;7388
                                                    P2_P2_P3_CodeFetch <= #1 1'b0; $display(";A 7389");		//(= P2_P2_P3_CodeFetch    0b0)) ;7389
                                                    P2_P2_P3_State2 = 4'sb0110; $display(";A 7390");		//(= P2_P2_P3_State2    0b0110)) ;7390
                                                end
                                                else begin
                                                    $display(";A 7384");		//(= (bv-comp P2_P2_P3_StateBS16  0b0)   0b0)) ;7384
                                                end
                                                P2_P2_P3_More = 1'b0; $display(";A 7391");		//(= P2_P2_P3_More    0b0)) ;7391
                                                P2_P2_P3_Flush = 1'b0; $display(";A 7392");		//(= P2_P2_P3_Flush    0b0)) ;7392
                                                P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7393");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;7393
                                                P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 7394");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;7394
                                            end
                                            else begin
                                                $display(";A 7381");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7381
                                            end
                                        end
                                        else begin
                                            $display(";A 7378");		//(= (bv-or (bv-comp P2_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P3_State  0b00000000000000000000000000000100))   0b0)) ;7378
                                        end
                                    end
                                    else begin
                                        $display(";A 7366");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;7366
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7395");		//(= P2_P2_P3_Flush    0b0)) ;7395
                                        P2_P2_P3_More = 1'b1; $display(";A 7396");		//(= P2_P2_P3_More    0b1)) ;7396
                                    end
                                end
                            8'b11100100 :
                                begin
                                    $display(";A 7397");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b11100100)) ;7397
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 7398");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;7398
                                        P2_P2_P3_rEIP <= #1 (P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 7400");		//(= P2_P2_P3_rEIP    (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;7400
                                        P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7401");		//(= P2_P2_P3_RequestPending    0b1)) ;7401
                                        P2_P2_P3_ReadRequest <= #1 1'b1; $display(";A 7402");		//(= P2_P2_P3_ReadRequest    0b1)) ;7402
                                        P2_P2_P3_MemoryFetch <= #1 1'b0; $display(";A 7403");		//(= P2_P2_P3_MemoryFetch    0b0)) ;7403
                                        P2_P2_P3_CodeFetch <= #1 1'b0; $display(";A 7404");		//(= P2_P2_P3_CodeFetch    0b0)) ;7404
                                        if ((P2_P2_P3_READY_n == 1'b0)) begin
                                            $display(";A 7405");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7405
                                            P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7407");		//(= P2_P2_P3_RequestPending    0b0)) ;7407
                                            P2_P2_P3_EAX <= #1 P2_P2_P3_Datai; $display(";A 7408");		//(= P2_P2_P3_EAX    P2_P2_P3_Datai )) ;7408
                                            P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7409");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;7409
                                            P2_P2_P3_InstQueueRd_Addr = (P2_P2_P3_InstQueueRd_Addr + 5'b00010); $display(";A 7410");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-add P2_P2_P3_InstQueueRd_Addr  0b00010))) ;7410
                                            P2_P2_P3_Flush = 1'b0; $display(";A 7411");		//(= P2_P2_P3_Flush    0b0)) ;7411
                                            P2_P2_P3_More = 1'b0; $display(";A 7412");		//(= P2_P2_P3_More    0b0)) ;7412
                                        end
                                        else begin
                                            $display(";A 7406");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7406
                                        end
                                    end
                                    else begin
                                        $display(";A 7399");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;7399
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7413");		//(= P2_P2_P3_Flush    0b0)) ;7413
                                        P2_P2_P3_More = 1'b1; $display(";A 7414");		//(= P2_P2_P3_More    0b1)) ;7414
                                    end
                                end
                            8'b11100110 :
                                begin
                                    $display(";A 7415");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b11100110)) ;7415
                                    if (((P2_P2_P3_InstQueueWr_Addr - P2_P2_P3_InstQueueRd_Addr) >= 32'b00000000000000000000000000000010)) begin
                                        $display(";A 7416");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b1)) ;7416
                                        P2_P2_P3_rEIP <= #1 (P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001); $display(";A 7418");		//(= P2_P2_P3_rEIP    (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001))) ;7418
                                        P2_P2_P3_RequestPending <= #1 1'b1; $display(";A 7419");		//(= P2_P2_P3_RequestPending    0b1)) ;7419
                                        P2_P2_P3_ReadRequest <= #1 1'b0; $display(";A 7420");		//(= P2_P2_P3_ReadRequest    0b0)) ;7420
                                        P2_P2_P3_MemoryFetch <= #1 1'b0; $display(";A 7421");		//(= P2_P2_P3_MemoryFetch    0b0)) ;7421
                                        P2_P2_P3_CodeFetch <= #1 1'b0; $display(";A 7422");		//(= P2_P2_P3_CodeFetch    0b0)) ;7422
                                        if (((P2_P2_P3_State == 32'b00000000000000000000000000000010) | (P2_P2_P3_State == 32'b00000000000000000000000000000100))) begin
                                            $display(";A 7423");		//(= (bv-or (bv-comp P2_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P3_State  0b00000000000000000000000000000100))   0b1)) ;7423
                                            P2_P2_P3_fWord = (P2_P2_P3_EAX % 32'b00000000000000010000000000000000); $display(";A 7425");		//(= P2_P2_P3_fWord    (bv-smod P2_P2_P3_EAX  0b00000000000000010000000000000000))) ;7425
                                            P2_P2_P3_Datao <= #1 P2_P2_P3_fWord; $display(";A 7426");		//(= P2_P2_P3_Datao    P2_P2_P3_fWord )) ;7426
                                            if ((P2_P2_P3_READY_n == 1'b0)) begin
                                                $display(";A 7427");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7427
                                                P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7429");		//(= P2_P2_P3_RequestPending    0b0)) ;7429
                                                P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7430");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;7430
                                                P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 7431");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;7431
                                                P2_P2_P3_Flush = 1'b0; $display(";A 7432");		//(= P2_P2_P3_Flush    0b0)) ;7432
                                                P2_P2_P3_More = 1'b0; $display(";A 7433");		//(= P2_P2_P3_More    0b0)) ;7433
                                            end
                                            else begin
                                                $display(";A 7428");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7428
                                            end
                                        end
                                        else begin
                                            $display(";A 7424");		//(= (bv-or (bv-comp P2_P2_P3_State  0b00000000000000000000000000000010) (bv-comp P2_P2_P3_State  0b00000000000000000000000000000100))   0b0)) ;7424
                                        end
                                    end
                                    else begin
                                        $display(";A 7417");		//(= (bool-to-bv (bv-ge (bv-sub P2_P2_P3_InstQueueWr_Addr  P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000010))   0b0)) ;7417
                                        P2_P2_P3_Flush = 1'b0; $display(";A 7434");		//(= P2_P2_P3_Flush    0b0)) ;7434
                                        P2_P2_P3_More = 1'b1; $display(";A 7435");		//(= P2_P2_P3_More    0b1)) ;7435
                                    end
                                end
                            8'b00000100 :
                                begin
                                    $display(";A 7436");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b00000100)) ;7436
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7437");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7437
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7438");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7438
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7439");		//(= P2_P2_P3_Flush    0b0)) ;7439
                                    P2_P2_P3_More = 1'b0; $display(";A 7440");		//(= P2_P2_P3_More    0b0)) ;7440
                                end
                            8'b00000101 :
                                begin
                                    $display(";A 7441");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b00000101)) ;7441
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7442");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7442
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7443");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7443
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7444");		//(= P2_P2_P3_Flush    0b0)) ;7444
                                    P2_P2_P3_More = 1'b0; $display(";A 7445");		//(= P2_P2_P3_More    0b0)) ;7445
                                end
                            8'b11010000 :
                                begin
                                    $display(";A 7446");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b11010000)) ;7446
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7447");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;7447
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 7448");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;7448
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7449");		//(= P2_P2_P3_Flush    0b0)) ;7449
                                    P2_P2_P3_More = 1'b0; $display(";A 7450");		//(= P2_P2_P3_More    0b0)) ;7450
                                end
                            8'b11000000 :
                                begin
                                    $display(";A 7451");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b11000000)) ;7451
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000010); $display(";A 7452");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000010))) ;7452
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000010) % 32'b00000000000000000000000000010000); $display(";A 7453");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000010) 0b00000000000000000000000000010000))) ;7453
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7454");		//(= P2_P2_P3_Flush    0b0)) ;7454
                                    P2_P2_P3_More = 1'b0; $display(";A 7455");		//(= P2_P2_P3_More    0b0)) ;7455
                                end
                            8'b01000000 :
                                begin
                                    $display(";A 7456");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b01000000)) ;7456
                                    P2_P2_P3_EAX <= #1 (P2_P2_P3_EAX + 32'sb00000000000000000000000000000001); $display(";A 7457");		//(= P2_P2_P3_EAX    (bv-add P2_P2_P3_EAX  0b00000000000000000000000000000001))) ;7457
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7458");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7458
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7459");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7459
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7460");		//(= P2_P2_P3_Flush    0b0)) ;7460
                                    P2_P2_P3_More = 1'b0; $display(";A 7461");		//(= P2_P2_P3_More    0b0)) ;7461
                                end
                            8'b01000011 :
                                begin
                                    $display(";A 7462");		//(= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr )   0b01000011)) ;7462
                                    P2_P2_P3_EBX <= #1 (P2_P2_P3_EBX + 32'sb00000000000000000000000000000001); $display(";A 7463");		//(= P2_P2_P3_EBX    (bv-add P2_P2_P3_EBX  0b00000000000000000000000000000001))) ;7463
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7464");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7464
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7465");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7465
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7466");		//(= P2_P2_P3_Flush    0b0)) ;7466
                                    P2_P2_P3_More = 1'b0; $display(";A 7467");		//(= P2_P2_P3_More    0b0)) ;7467
                                end
                            default:
                                begin
                                    $display(";A 7468");		//(= (and (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b10010000) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b01100110) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b11101011) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b11101001) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b11101010) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b10110000) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b10111000) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b10111011) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b10001011) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b10001001) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b11100100) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b11100110) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b00000100) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b00000101) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b11010000) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b11000000) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b01000000) (/= ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ) 0b01000011))   true)) ;7468
                                    P2_P2_P3_InstAddrPointer = (P2_P2_P3_InstAddrPointer + 32'sb00000000000000000000000000000001); $display(";A 7469");		//(= P2_P2_P3_InstAddrPointer    (bv-add P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000001))) ;7469
                                    P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7470");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7470
                                    P2_P2_P3_Flush = 1'b0; $display(";A 7471");		//(= P2_P2_P3_Flush    0b0)) ;7471
                                    P2_P2_P3_More = 1'b0; $display(";A 7472");		//(= P2_P2_P3_More    0b0)) ;7472
                                end
                        endcase
                        if (((~(P2_P2_P3_InstQueueRd_Addr < P2_P2_P3_InstQueueWr_Addr)) | ((((32'b00000000000000000000000000001111 - P2_P2_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000100) | P2_P2_P3_Flush) | P2_P2_P3_More))) begin
                            $display(";A 7473");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P2_P3_InstQueueRd_Addr  P2_P2_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P2_P3_Flush ) P2_P2_P3_More ))   0b1)) ;7473
                            P2_P2_P3_State2 = 4'sb0111; $display(";A 7475");		//(= P2_P2_P3_State2    0b0111)) ;7475
                        end
                        else begin
                            $display(";A 7474");		//(= (bv-or (bv-not (bool-to-bv (bv-lt P2_P2_P3_InstQueueRd_Addr  P2_P2_P3_InstQueueWr_Addr ))) (bv-or (bv-or (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000100)) P2_P2_P3_Flush ) P2_P2_P3_More ))   0b0)) ;7474
                        end
                    end
                4'b0110 :
                    begin
                        $display(";A 7476");		//(= P2_P2_P3_State2    0b0110)) ;7476
                        P2_P2_P3_Datao <= #1 ((P2_P2_P3_uWord * 32'b00000000000000010000000000000000) + P2_P2_P3_lWord); $display(";A 7477");		//(= P2_P2_P3_Datao    (bv-add (bv-mul P2_P2_P3_uWord  0b00000000000000010000000000000000) P2_P2_P3_lWord ))) ;7477
                        if ((P2_P2_P3_READY_n == 1'b0)) begin
                            $display(";A 7478");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b1)) ;7478
                            P2_P2_P3_RequestPending <= #1 1'b0; $display(";A 7480");		//(= P2_P2_P3_RequestPending    0b0)) ;7480
                            P2_P2_P3_State2 = 4'sb0101; $display(";A 7481");		//(= P2_P2_P3_State2    0b0101)) ;7481
                        end
                        else begin
                            $display(";A 7479");		//(= (bv-comp P2_P2_P3_READY_n  0b0)   0b0)) ;7479
                        end
                    end
                4'b0111 :
                    begin
                        $display(";A 7482");		//(= P2_P2_P3_State2    0b0111)) ;7482
                        if (P2_P2_P3_Flush) begin
                            $display(";A 7483");		//(= P2_P2_P3_Flush    0b1)) ;7483
                            P2_P2_P3_InstQueueRd_Addr = 5'sb00001; $display(";A 7485");		//(= P2_P2_P3_InstQueueRd_Addr    0b00001)) ;7485
                            P2_P2_P3_InstQueueWr_Addr = 5'sb00001; $display(";A 7486");		//(= P2_P2_P3_InstQueueWr_Addr    0b00001)) ;7486
                            if ((P2_P2_P3_InstAddrPointer < 32'sb00000000000000000000000000000000)) begin
                                $display(";A 7487");		//(= (bool-to-bv (bv-slt P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b1)) ;7487
                                P2_P2_P3_fWord = (-P2_P2_P3_InstAddrPointer); $display(";A 7489");		//(= P2_P2_P3_fWord    (bv-neg P2_P2_P3_InstAddrPointer ))) ;7489
                            end
                            else begin
                                $display(";A 7488");		//(= (bool-to-bv (bv-slt P2_P2_P3_InstAddrPointer  0b00000000000000000000000000000000))   0b0)) ;7488
                                P2_P2_P3_fWord = P2_P2_P3_InstAddrPointer; $display(";A 7490");		//(= P2_P2_P3_fWord    P2_P2_P3_InstAddrPointer )) ;7490
                            end
                            if (((P2_P2_P3_fWord % 32'sb00000000000000000000000000000010) == 32'sb00000000000000000000000000000001)) begin
                                $display(";A 7491");		//(= (bv-comp (bv-smod P2_P2_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b1)) ;7491
                                P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + (P2_P2_P3_fWord % 32'b00000000000000000000000000000100)) % 32'b00000000000000000000000000010000); $display(";A 7493");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  (bv-smod P2_P2_P3_fWord  0b00000000000000000000000000000100)) 0b00000000000000000000000000010000))) ;7493
                            end
                            else begin
                                $display(";A 7492");		//(= (bv-comp (bv-smod P2_P2_P3_fWord  0b00000000000000000000000000000010) 0b00000000000000000000000000000001)   0b0)) ;7492
                            end
                        end
                        else begin
                            $display(";A 7484");		//(= P2_P2_P3_Flush    0b0)) ;7484
                        end
                        if (((32'b00000000000000000000000000001111 - P2_P2_P3_InstQueueRd_Addr) < 32'b00000000000000000000000000000011)) begin
                            $display(";A 7494");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b1)) ;7494
                            P2_P2_P3_State2 = 4'sb1000; $display(";A 7496");		//(= P2_P2_P3_State2    0b1000)) ;7496
                            P2_P2_P3_InstQueueWr_Addr = 5'sb00000; $display(";A 7497");		//(= P2_P2_P3_InstQueueWr_Addr    0b00000)) ;7497
                        end
                        else begin
                            $display(";A 7495");		//(= (bool-to-bv (bv-lt (bv-sub 0b00000000000000000000000000001111 P2_P2_P3_InstQueueRd_Addr ) 0b00000000000000000000000000000011))   0b0)) ;7495
                            P2_P2_P3_State2 = 4'sb1001; $display(";A 7498");		//(= P2_P2_P3_State2    0b1001)) ;7498
                        end
                    end
                4'b1000 :
                    begin
                        $display(";A 7499");		//(= P2_P2_P3_State2    0b1000)) ;7499
                        if ((P2_P2_P3_InstQueueRd_Addr <= 32'b00000000000000000000000000001111)) begin
                            $display(";A 7500");		//(= (bool-to-bv (bv-le P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b1)) ;7500
                            P2_P2_P3_InstQueue[P2_P2_P3_InstQueueWr_Addr] = P2_P2_P3_InstQueue[P2_P2_P3_InstQueueRd_Addr]; $display(";A 7502");		//(= P2_P2_P3_InstQueue    ( P2_P2_P3_InstQueue P2_P2_P3_InstQueueRd_Addr ))) ;7502
                            P2_P2_P3_InstQueueRd_Addr = ((P2_P2_P3_InstQueueRd_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7503");		//(= P2_P2_P3_InstQueueRd_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7503
                            P2_P2_P3_InstQueueWr_Addr = ((P2_P2_P3_InstQueueWr_Addr + 32'b00000000000000000000000000000001) % 32'b00000000000000000000000000010000); $display(";A 7504");		//(= P2_P2_P3_InstQueueWr_Addr    (bv-smod (bv-add P2_P2_P3_InstQueueWr_Addr  0b00000000000000000000000000000001) 0b00000000000000000000000000010000))) ;7504
                            P2_P2_P3_State2 = 4'sb1000; $display(";A 7505");		//(= P2_P2_P3_State2    0b1000)) ;7505
                        end
                        else begin
                            $display(";A 7501");		//(= (bool-to-bv (bv-le P2_P2_P3_InstQueueRd_Addr  0b00000000000000000000000000001111))   0b0)) ;7501
                            P2_P2_P3_InstQueueRd_Addr = 5'sb00000; $display(";A 7506");		//(= P2_P2_P3_InstQueueRd_Addr    0b00000)) ;7506
                            P2_P2_P3_State2 = 4'sb1001; $display(";A 7507");		//(= P2_P2_P3_State2    0b1001)) ;7507
                        end
                    end
                4'b1001 :
                    begin
                        $display(";A 7508");		//(= P2_P2_P3_State2    0b1001)) ;7508
                        P2_P2_P3_rEIP <= #1 P2_P2_P3_PhyAddrPointer; $display(";A 7509");		//(= P2_P2_P3_rEIP    P2_P2_P3_PhyAddrPointer )) ;7509
                        P2_P2_P3_State2 = 4'sb0001; $display(";A 7510");		//(= P2_P2_P3_State2    0b0001)) ;7510
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:11487
    always @(posedge P2_P2_P3_RESET or posedge P2_P2_P3_CLOCK) begin
        if ((P2_P2_P3_RESET == 1'b1)) begin
            $display(";A 7511");		//(= (bv-comp P2_P2_P3_RESET  0b1)   0b1)) ;7511
            P2_P2_P3_ByteEnable <= #1 4'b0000; $display(";A 7513");		//(= P2_P2_P3_ByteEnable    0b0000)) ;7513
            P2_P2_P3_NonAligned <= #1 1'b0; $display(";A 7514");		//(= P2_P2_P3_NonAligned    0b0)) ;7514
        end
        else begin
            $display(";A 7512");		//(= (bv-comp P2_P2_P3_RESET  0b1)   0b0)) ;7512
            case (P2_P2_P3_DataWidth)
                32'sb00000000000000000000000000000000 :
                    begin
                        $display(";A 7515");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000000)) ;7515
                        case ((P2_P2_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 7516");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;7516
                                    P2_P2_P3_ByteEnable <= #1 4'b1110; $display(";A 7517");		//(= P2_P2_P3_ByteEnable    0b1110)) ;7517
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 7518");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;7518
                                    P2_P2_P3_ByteEnable <= #1 4'b1101; $display(";A 7519");		//(= P2_P2_P3_ByteEnable    0b1101)) ;7519
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 7520");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;7520
                                    P2_P2_P3_ByteEnable <= #1 4'b1011; $display(";A 7521");		//(= P2_P2_P3_ByteEnable    0b1011)) ;7521
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 7522");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;7522
                                    P2_P2_P3_ByteEnable <= #1 4'b0111; $display(";A 7523");		//(= P2_P2_P3_ByteEnable    0b0111)) ;7523
                                end
                            default:
                                begin
                                    $display(";A 7524");		//(= (and (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;7524
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000001 :
                    begin
                        $display(";A 7525");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000001)) ;7525
                        case ((P2_P2_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 7526");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;7526
                                    P2_P2_P3_ByteEnable <= #1 4'b1100; $display(";A 7527");		//(= P2_P2_P3_ByteEnable    0b1100)) ;7527
                                    P2_P2_P3_NonAligned <= #1 1'b0; $display(";A 7528");		//(= P2_P2_P3_NonAligned    0b0)) ;7528
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 7529");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;7529
                                    P2_P2_P3_ByteEnable <= #1 4'b1001; $display(";A 7530");		//(= P2_P2_P3_ByteEnable    0b1001)) ;7530
                                    P2_P2_P3_NonAligned <= #1 1'b0; $display(";A 7531");		//(= P2_P2_P3_NonAligned    0b0)) ;7531
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 7532");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;7532
                                    P2_P2_P3_ByteEnable <= #1 4'b0011; $display(";A 7533");		//(= P2_P2_P3_ByteEnable    0b0011)) ;7533
                                    P2_P2_P3_NonAligned <= #1 1'b0; $display(";A 7534");		//(= P2_P2_P3_NonAligned    0b0)) ;7534
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 7535");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;7535
                                    P2_P2_P3_ByteEnable <= #1 4'b0111; $display(";A 7536");		//(= P2_P2_P3_ByteEnable    0b0111)) ;7536
                                    P2_P2_P3_NonAligned <= #1 1'b1; $display(";A 7537");		//(= P2_P2_P3_NonAligned    0b1)) ;7537
                                end
                            default:
                                begin
                                    $display(";A 7538");		//(= (and (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;7538
                                    begin
                                    end
                                end
                        endcase
                    end
                32'sb00000000000000000000000000000010 :
                    begin
                        $display(";A 7539");		//(= P2_P2_P3_DataWidth    0b00000000000000000000000000000010)) ;7539
                        case ((P2_P2_P3_rEIP % 32'sb00000000000000000000000000000100))
                            32'sb00000000000000000000000000000000 :
                                begin
                                    $display(";A 7540");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000000)) ;7540
                                    P2_P2_P3_ByteEnable <= #1 4'b0000; $display(";A 7541");		//(= P2_P2_P3_ByteEnable    0b0000)) ;7541
                                    P2_P2_P3_NonAligned <= #1 1'b0; $display(";A 7542");		//(= P2_P2_P3_NonAligned    0b0)) ;7542
                                end
                            32'sb00000000000000000000000000000001 :
                                begin
                                    $display(";A 7543");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000001)) ;7543
                                    P2_P2_P3_ByteEnable <= #1 4'b0001; $display(";A 7544");		//(= P2_P2_P3_ByteEnable    0b0001)) ;7544
                                    P2_P2_P3_NonAligned <= #1 1'b1; $display(";A 7545");		//(= P2_P2_P3_NonAligned    0b1)) ;7545
                                end
                            32'sb00000000000000000000000000000010 :
                                begin
                                    $display(";A 7546");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000010)) ;7546
                                    P2_P2_P3_NonAligned <= #1 1'b1; $display(";A 7547");		//(= P2_P2_P3_NonAligned    0b1)) ;7547
                                    P2_P2_P3_ByteEnable <= #1 4'b0011; $display(";A 7548");		//(= P2_P2_P3_ByteEnable    0b0011)) ;7548
                                end
                            32'sb00000000000000000000000000000011 :
                                begin
                                    $display(";A 7549");		//(= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100)   0b00000000000000000000000000000011)) ;7549
                                    P2_P2_P3_NonAligned <= #1 1'b1; $display(";A 7550");		//(= P2_P2_P3_NonAligned    0b1)) ;7550
                                    P2_P2_P3_ByteEnable <= #1 4'b0111; $display(";A 7551");		//(= P2_P2_P3_ByteEnable    0b0111)) ;7551
                                end
                            default:
                                begin
                                    $display(";A 7552");		//(= (and (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000000) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000001) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000010) (/= (bv-smod P2_P2_P3_rEIP  0b00000000000000000000000000000100) 0b00000000000000000000000000000011))   true)) ;7552
                                    begin
                                    end
                                end
                        endcase
                    end
                default:
                    begin
                        $display(";A 7553");		//(= (and (/= P2_P2_P3_DataWidth  0b00000000000000000000000000000000) (/= P2_P2_P3_DataWidth  0b00000000000000000000000000000001) (/= P2_P2_P3_DataWidth  0b00000000000000000000000000000010))   true)) ;7553
                        begin
                        end
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:11604
    always @(posedge P2_P3_reset or posedge P2_P3_clock) begin
        if ((P2_P3_reset == 1'b1)) begin
            P2_P3_MAR = 20'sb00000000000000000000; $display(";A 7556");		//(= P2_P3_MAR    0b00000000000000000000)) ;7556
            P2_P3_MBR = 32'sb00000000000000000000000000000000; $display(";A 7557");		//(= P2_P3_MBR    0b00000000000000000000000000000000)) ;7557
            P2_P3_IR = 32'sb00000000000000000000000000000000; $display(";A 7558");		//(= P2_P3_IR    0b00000000000000000000000000000000)) ;7558
            P2_P3_d = 32'sb00000000000000000000000000000000; $display(";A 7559");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7559
            P2_P3_r = 32'sb00000000000000000000000000000000; $display(";A 7560");		//(= P2_P3_r    0b00000000000000000000000000000000)) ;7560
            P2_P3_m = 32'sb00000000000000000000000000000000; $display(";A 7561");		//(= P2_P3_m    0b00000000000000000000000000000000)) ;7561
            P2_P3_s = 2'sb00; $display(";A 7562");		//(= P2_P3_s    0b00)) ;7562
            P2_P3_temp = 32'sb00000000000000000000000000000000; $display(";A 7563");		//(= P2_P3_temp    0b00000000000000000000000000000000)) ;7563
            P2_P3_mf = 2'sb00; $display(";A 7564");		//(= P2_P3_mf    0b00)) ;7564
            P2_P3_df = 3'sb000; $display(";A 7565");		//(= P2_P3_df    0b000)) ;7565
            P2_P3_ff = 4'sb0000; $display(";A 7566");		//(= P2_P3_ff    0b0000)) ;7566
            P2_P3_cf = 1'sb0; $display(";A 7567");		//(= P2_P3_cf    0b0)) ;7567
            P2_P3_tail = 20'sb00000000000000000000; $display(";A 7568");		//(= P2_P3_tail    0b00000000000000000000)) ;7568
            P2_P3_B = 1'b0; $display(";A 7569");		//(= P2_P3_B    0b0)) ;7569
            P2_P3_reg0 = 32'sb00000000000000000000000000000000; $display(";A 7570");		//(= P2_P3_reg0    0b00000000000000000000000000000000)) ;7570
            P2_P3_reg1 = 32'sb00000000000000000000000000000000; $display(";A 7571");		//(= P2_P3_reg1    0b00000000000000000000000000000000)) ;7571
            P2_P3_reg2 = 32'sb00000000000000000000000000000000; $display(";A 7572");		//(= P2_P3_reg2    0b00000000000000000000000000000000)) ;7572
            P2_P3_reg3 = 32'sb00000000000000000000000000000000; $display(";A 7573");		//(= P2_P3_reg3    0b00000000000000000000000000000000)) ;7573
            P2_P3_addr <= #1 20'sb00000000000000000000; $display(";A 7574");		//(= P2_P3_addr    0b00000000000000000000)) ;7574
            P2_P3_rd <= #1 1'b0; $display(";A 7575");		//(= P2_P3_rd    0b0)) ;7575
            P2_P3_wr <= #1 1'b0; $display(";A 7576");		//(= P2_P3_wr    0b0)) ;7576
            P2_P3_datao <= #1 32'sb00000000000000000000000000000000; $display(";A 7577");		//(= P2_P3_datao    0b00000000000000000000000000000000)) ;7577
            P2_P3_state = 1'sb0; $display(";A 7578");		//(= P2_P3_state    0b0)) ;7578
        end
        else begin
            P2_P3_rd <= #1 1'b0; $display(";A 7579");		//(= P2_P3_rd    0b0)) ;7579
            P2_P3_wr <= #1 1'b0; $display(";A 7580");		//(= P2_P3_wr    0b0)) ;7580
            case (P2_P3_state)
                1'b0 :
                    begin
                        $display(";A 7581");		//(= P2_P3_state    0b0)) ;7581
                        P2_P3_MAR = (P2_P3_reg3 % 32'b00000000000100000000000000000000); $display(";A 7582");		//(= P2_P3_MAR    (bv-smod P2_P3_reg3  0b00000000000100000000000000000000))) ;7582
                        P2_P3_addr <= #1 P2_P3_MAR; $display(";A 7583");		//(= P2_P3_addr    P2_P3_MAR )) ;7583
                        P2_P3_rd <= #1 1'b1; $display(";A 7584");		//(= P2_P3_rd    0b1)) ;7584
                        P2_P3_MBR = P2_P3_datai; $display(";A 7585");		//(= P2_P3_MBR    P2_P3_datai )) ;7585
                        P2_P3_IR = P2_P3_MBR; $display(";A 7586");		//(= P2_P3_IR    P2_P3_MBR )) ;7586
                        P2_P3_state = 1'sb1; $display(";A 7587");		//(= P2_P3_state    0b1)) ;7587
                    end
                1'b1 :
                    begin
                        $display(";A 7588");		//(= P2_P3_state    0b1)) ;7588
                        if ((P2_P3_IR < 32'sb00000000000000000000000000000000)) begin
                            $display(";A 7589");		//(= (bool-to-bv (bv-slt P2_P3_IR  0b00000000000000000000000000000000))   0b1)) ;7589
                            P2_P3_IR = (-P2_P3_IR); $display(";A 7591");		//(= P2_P3_IR    (bv-neg P2_P3_IR ))) ;7591
                        end
                        else begin
                            $display(";A 7590");		//(= (bool-to-bv (bv-slt P2_P3_IR  0b00000000000000000000000000000000))   0b0)) ;7590
                        end
                        P2_P3_mf = ((P2_P3_IR / 32'b00001000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 7592");		//(= P2_P3_mf    (bv-smod (bv-sdiv P2_P3_IR  0b00001000000000000000000000000000) 0b00000000000000000000000000000100))) ;7592
                        P2_P3_df = ((P2_P3_IR / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000000001000); $display(";A 7593");		//(= P2_P3_df    (bv-smod (bv-sdiv P2_P3_IR  0b00000001000000000000000000000000) 0b00000000000000000000000000001000))) ;7593
                        P2_P3_ff = ((P2_P3_IR / 32'b00000000000010000000000000000000) % 32'b00000000000000000000000000010000); $display(";A 7594");		//(= P2_P3_ff    (bv-smod (bv-sdiv P2_P3_IR  0b00000000000010000000000000000000) 0b00000000000000000000000000010000))) ;7594
                        P2_P3_cf = ((P2_P3_IR / 32'b00000000100000000000000000000000) % 32'b00000000000000000000000000000010); $display(";A 7595");		//(= P2_P3_cf    (bv-smod (bv-sdiv P2_P3_IR  0b00000000100000000000000000000000) 0b00000000000000000000000000000010))) ;7595
                        P2_P3_tail = (P2_P3_IR % 32'b00000000000100000000000000000000); $display(";A 7596");		//(= P2_P3_tail    (bv-smod P2_P3_IR  0b00000000000100000000000000000000))) ;7596
                        P2_P3_reg3 = ((P2_P3_reg3 % 32'b00100000000000000000000000000000) + 32'b00000000000000000000000000001000); $display(";A 7597");		//(= P2_P3_reg3    (bv-add (bv-smod P2_P3_reg3  0b00100000000000000000000000000000) 0b00000000000000000000000000001000))) ;7597
                        P2_P3_s = ((P2_P3_IR / 32'b00100000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 7598");		//(= P2_P3_s    (bv-smod (bv-sdiv P2_P3_IR  0b00100000000000000000000000000000) 0b00000000000000000000000000000100))) ;7598
                        case (P2_P3_s)
                            2'b00 :
                                begin
                                    $display(";A 7599");		//(= P2_P3_s    0b00)) ;7599
                                    P2_P3_r = P2_P3_reg0; $display(";A 7600");		//(= P2_P3_r    P2_P3_reg0 )) ;7600
                                end
                            2'b01 :
                                begin
                                    $display(";A 7601");		//(= P2_P3_s    0b01)) ;7601
                                    P2_P3_r = P2_P3_reg1; $display(";A 7602");		//(= P2_P3_r    P2_P3_reg1 )) ;7602
                                end
                            2'b10 :
                                begin
                                    $display(";A 7603");		//(= P2_P3_s    0b10)) ;7603
                                    P2_P3_r = P2_P3_reg2; $display(";A 7604");		//(= P2_P3_r    P2_P3_reg2 )) ;7604
                                end
                            2'b11 :
                                begin
                                    $display(";A 7605");		//(= P2_P3_s    0b11)) ;7605
                                    P2_P3_r = P2_P3_reg3; $display(";A 7606");		//(= P2_P3_r    P2_P3_reg3 )) ;7606
                                end
                        endcase
                        case (P2_P3_cf)
                            1'b1 :
                                begin
                                    $display(";A 7607");		//(= P2_P3_cf    0b1)) ;7607
                                    case (P2_P3_mf)
                                        2'b00 :
                                            begin
                                                $display(";A 7608");		//(= P2_P3_mf    0b00)) ;7608
                                                P2_P3_m = P2_P3_tail; $display(";A 7609");		//(= P2_P3_m    P2_P3_tail )) ;7609
                                            end
                                        2'b01 :
                                            begin
                                                $display(";A 7610");		//(= P2_P3_mf    0b01)) ;7610
                                                P2_P3_m = P2_P3_datai; $display(";A 7611");		//(= P2_P3_m    P2_P3_datai )) ;7611
                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7612");		//(= P2_P3_addr    P2_P3_tail )) ;7612
                                                P2_P3_rd <= #1 1'b1; $display(";A 7613");		//(= P2_P3_rd    0b1)) ;7613
                                            end
                                        2'b10 :
                                            begin
                                                $display(";A 7614");		//(= P2_P3_mf    0b10)) ;7614
                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7615");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7615
                                                P2_P3_rd <= #1 1'b1; $display(";A 7616");		//(= P2_P3_rd    0b1)) ;7616
                                                P2_P3_m = P2_P3_datai; $display(";A 7617");		//(= P2_P3_m    P2_P3_datai )) ;7617
                                            end
                                        2'b11 :
                                            begin
                                                $display(";A 7618");		//(= P2_P3_mf    0b11)) ;7618
                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7619");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7619
                                                P2_P3_rd <= #1 1'b1; $display(";A 7620");		//(= P2_P3_rd    0b1)) ;7620
                                                P2_P3_m = P2_P3_datai; $display(";A 7621");		//(= P2_P3_m    P2_P3_datai )) ;7621
                                            end
                                    endcase
                                    case (P2_P3_ff)
                                        4'b0000 :
                                            begin
                                                $display(";A 7622");		//(= P2_P3_ff    0b0000)) ;7622
                                                if ((P2_P3_r < P2_P3_m)) begin
                                                    $display(";A 7623");		//(= (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))   0b1)) ;7623
                                                    P2_P3_B = 1'b1; $display(";A 7625");		//(= P2_P3_B    0b1)) ;7625
                                                end
                                                else begin
                                                    $display(";A 7624");		//(= (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))   0b0)) ;7624
                                                    P2_P3_B = 1'b0; $display(";A 7626");		//(= P2_P3_B    0b0)) ;7626
                                                end
                                            end
                                        4'b0001 :
                                            begin
                                                $display(";A 7627");		//(= P2_P3_ff    0b0001)) ;7627
                                                if ((~(P2_P3_r < P2_P3_m))) begin
                                                    $display(";A 7628");		//(= (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )))   0b1)) ;7628
                                                    P2_P3_B = 1'b1; $display(";A 7630");		//(= P2_P3_B    0b1)) ;7630
                                                end
                                                else begin
                                                    $display(";A 7629");		//(= (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )))   0b0)) ;7629
                                                    P2_P3_B = 1'b0; $display(";A 7631");		//(= P2_P3_B    0b0)) ;7631
                                                end
                                            end
                                        4'b0010 :
                                            begin
                                                $display(";A 7632");		//(= P2_P3_ff    0b0010)) ;7632
                                                if ((P2_P3_r == P2_P3_m)) begin
                                                    $display(";A 7633");		//(= (bv-comp P2_P3_r  P2_P3_m )   0b1)) ;7633
                                                    P2_P3_B = 1'b1; $display(";A 7635");		//(= P2_P3_B    0b1)) ;7635
                                                end
                                                else begin
                                                    $display(";A 7634");		//(= (bv-comp P2_P3_r  P2_P3_m )   0b0)) ;7634
                                                    P2_P3_B = 1'b0; $display(";A 7636");		//(= P2_P3_B    0b0)) ;7636
                                                end
                                            end
                                        4'b0011 :
                                            begin
                                                $display(";A 7637");		//(= P2_P3_ff    0b0011)) ;7637
                                                if ((~(P2_P3_r == P2_P3_m))) begin
                                                    $display(";A 7638");		//(= (bv-not (bv-comp P2_P3_r  P2_P3_m ))   0b1)) ;7638
                                                    P2_P3_B = 1'b1; $display(";A 7640");		//(= P2_P3_B    0b1)) ;7640
                                                end
                                                else begin
                                                    $display(";A 7639");		//(= (bv-not (bv-comp P2_P3_r  P2_P3_m ))   0b0)) ;7639
                                                    P2_P3_B = 1'b0; $display(";A 7641");		//(= P2_P3_B    0b0)) ;7641
                                                end
                                            end
                                        4'b0100 :
                                            begin
                                                $display(";A 7642");		//(= P2_P3_ff    0b0100)) ;7642
                                                if ((~(P2_P3_r > P2_P3_m))) begin
                                                    $display(";A 7643");		//(= (bv-not (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m )))   0b1)) ;7643
                                                    P2_P3_B = 1'b1; $display(";A 7645");		//(= P2_P3_B    0b1)) ;7645
                                                end
                                                else begin
                                                    $display(";A 7644");		//(= (bv-not (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m )))   0b0)) ;7644
                                                    P2_P3_B = 1'b0; $display(";A 7646");		//(= P2_P3_B    0b0)) ;7646
                                                end
                                            end
                                        4'b0101 :
                                            begin
                                                $display(";A 7647");		//(= P2_P3_ff    0b0101)) ;7647
                                                if ((P2_P3_r > P2_P3_m)) begin
                                                    $display(";A 7648");		//(= (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m ))   0b1)) ;7648
                                                    P2_P3_B = 1'b1; $display(";A 7650");		//(= P2_P3_B    0b1)) ;7650
                                                end
                                                else begin
                                                    $display(";A 7649");		//(= (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m ))   0b0)) ;7649
                                                    P2_P3_B = 1'b0; $display(";A 7651");		//(= P2_P3_B    0b0)) ;7651
                                                end
                                            end
                                        4'b0110 :
                                            begin
                                                $display(";A 7652");		//(= P2_P3_ff    0b0110)) ;7652
                                                if ((P2_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 7653");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b1)) ;7653
                                                    P2_P3_r = (P2_P3_r - 32'b00000000000000000000000000000000); $display(";A 7655");		//(= P2_P3_r    (bv-sub P2_P3_r  0b00000000000000000000000000000000))) ;7655
                                                end
                                                else begin
                                                    $display(";A 7654");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b0)) ;7654
                                                end
                                                if ((P2_P3_r < P2_P3_m)) begin
                                                    $display(";A 7656");		//(= (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))   0b1)) ;7656
                                                    P2_P3_B = 1'b1; $display(";A 7658");		//(= P2_P3_B    0b1)) ;7658
                                                end
                                                else begin
                                                    $display(";A 7657");		//(= (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))   0b0)) ;7657
                                                    P2_P3_B = 1'b0; $display(";A 7659");		//(= P2_P3_B    0b0)) ;7659
                                                end
                                            end
                                        4'b0111 :
                                            begin
                                                $display(";A 7660");		//(= P2_P3_ff    0b0111)) ;7660
                                                if ((P2_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 7661");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b1)) ;7661
                                                    P2_P3_r = (P2_P3_r - 32'b00000000000000000000000000000000); $display(";A 7663");		//(= P2_P3_r    (bv-sub P2_P3_r  0b00000000000000000000000000000000))) ;7663
                                                end
                                                else begin
                                                    $display(";A 7662");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b0)) ;7662
                                                end
                                                if ((~(P2_P3_r < P2_P3_m))) begin
                                                    $display(";A 7664");		//(= (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )))   0b1)) ;7664
                                                    P2_P3_B = 1'b1; $display(";A 7666");		//(= P2_P3_B    0b1)) ;7666
                                                end
                                                else begin
                                                    $display(";A 7665");		//(= (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )))   0b0)) ;7665
                                                    P2_P3_B = 1'b0; $display(";A 7667");		//(= P2_P3_B    0b0)) ;7667
                                                end
                                            end
                                        4'b1000 :
                                            begin
                                                $display(";A 7668");		//(= P2_P3_ff    0b1000)) ;7668
                                                if (((P2_P3_r < P2_P3_m) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7669");		//(= (bv-or (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b1)) ;7669
                                                    P2_P3_B = 1'b1; $display(";A 7671");		//(= P2_P3_B    0b1)) ;7671
                                                end
                                                else begin
                                                    $display(";A 7670");		//(= (bv-or (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b0)) ;7670
                                                    P2_P3_B = 1'b0; $display(";A 7672");		//(= P2_P3_B    0b0)) ;7672
                                                end
                                            end
                                        4'b1001 :
                                            begin
                                                $display(";A 7673");		//(= P2_P3_ff    0b1001)) ;7673
                                                if (((~(P2_P3_r < P2_P3_m)) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7674");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))) (bv-comp P2_P3_B  0b1))   0b1)) ;7674
                                                    P2_P3_B = 1'b1; $display(";A 7676");		//(= P2_P3_B    0b1)) ;7676
                                                end
                                                else begin
                                                    $display(";A 7675");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))) (bv-comp P2_P3_B  0b1))   0b0)) ;7675
                                                    P2_P3_B = 1'b0; $display(";A 7677");		//(= P2_P3_B    0b0)) ;7677
                                                end
                                            end
                                        4'b1010 :
                                            begin
                                                $display(";A 7678");		//(= P2_P3_ff    0b1010)) ;7678
                                                if (((P2_P3_r == P2_P3_m) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7679");		//(= (bv-or (bv-comp P2_P3_r  P2_P3_m ) (bv-comp P2_P3_B  0b1))   0b1)) ;7679
                                                    P2_P3_B = 1'b1; $display(";A 7681");		//(= P2_P3_B    0b1)) ;7681
                                                end
                                                else begin
                                                    $display(";A 7680");		//(= (bv-or (bv-comp P2_P3_r  P2_P3_m ) (bv-comp P2_P3_B  0b1))   0b0)) ;7680
                                                    P2_P3_B = 1'b0; $display(";A 7682");		//(= P2_P3_B    0b0)) ;7682
                                                end
                                            end
                                        4'b1011 :
                                            begin
                                                $display(";A 7683");		//(= P2_P3_ff    0b1011)) ;7683
                                                if (((~(P2_P3_r == P2_P3_m)) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7684");		//(= (bv-or (bv-not (bv-comp P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b1)) ;7684
                                                    P2_P3_B = 1'b1; $display(";A 7686");		//(= P2_P3_B    0b1)) ;7686
                                                end
                                                else begin
                                                    $display(";A 7685");		//(= (bv-or (bv-not (bv-comp P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b0)) ;7685
                                                    P2_P3_B = 1'b0; $display(";A 7687");		//(= P2_P3_B    0b0)) ;7687
                                                end
                                            end
                                        4'b1100 :
                                            begin
                                                $display(";A 7688");		//(= P2_P3_ff    0b1100)) ;7688
                                                if (((~(P2_P3_r > P2_P3_m)) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7689");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m ))) (bv-comp P2_P3_B  0b1))   0b1)) ;7689
                                                    P2_P3_B = 1'b1; $display(";A 7691");		//(= P2_P3_B    0b1)) ;7691
                                                end
                                                else begin
                                                    $display(";A 7690");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m ))) (bv-comp P2_P3_B  0b1))   0b0)) ;7690
                                                    P2_P3_B = 1'b0; $display(";A 7692");		//(= P2_P3_B    0b0)) ;7692
                                                end
                                            end
                                        4'b1101 :
                                            begin
                                                $display(";A 7693");		//(= P2_P3_ff    0b1101)) ;7693
                                                if (((P2_P3_r > P2_P3_m) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7694");		//(= (bv-or (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b1)) ;7694
                                                    P2_P3_B = 1'b1; $display(";A 7696");		//(= P2_P3_B    0b1)) ;7696
                                                end
                                                else begin
                                                    $display(";A 7695");		//(= (bv-or (bool-to-bv (bv-sgt P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b0)) ;7695
                                                    P2_P3_B = 1'b0; $display(";A 7697");		//(= P2_P3_B    0b0)) ;7697
                                                end
                                            end
                                        4'b1110 :
                                            begin
                                                $display(";A 7698");		//(= P2_P3_ff    0b1110)) ;7698
                                                if ((P2_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 7699");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b1)) ;7699
                                                    P2_P3_r = (P2_P3_r - 32'b00000000000000000000000000000000); $display(";A 7701");		//(= P2_P3_r    (bv-sub P2_P3_r  0b00000000000000000000000000000000))) ;7701
                                                end
                                                else begin
                                                    $display(";A 7700");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b0)) ;7700
                                                end
                                                if (((P2_P3_r < P2_P3_m) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7702");		//(= (bv-or (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b1)) ;7702
                                                    P2_P3_B = 1'b1; $display(";A 7704");		//(= P2_P3_B    0b1)) ;7704
                                                end
                                                else begin
                                                    $display(";A 7703");		//(= (bv-or (bool-to-bv (bv-slt P2_P3_r  P2_P3_m )) (bv-comp P2_P3_B  0b1))   0b0)) ;7703
                                                    P2_P3_B = 1'b0; $display(";A 7705");		//(= P2_P3_B    0b0)) ;7705
                                                end
                                            end
                                        4'b1111 :
                                            begin
                                                $display(";A 7706");		//(= P2_P3_ff    0b1111)) ;7706
                                                if ((P2_P3_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 7707");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b1)) ;7707
                                                    P2_P3_r = (P2_P3_r - 32'b00000000000000000000000000000000); $display(";A 7709");		//(= P2_P3_r    (bv-sub P2_P3_r  0b00000000000000000000000000000000))) ;7709
                                                end
                                                else begin
                                                    $display(";A 7708");		//(= (bool-to-bv (bv-gt P2_P3_r  0b11111111111111111111111111111111))   0b0)) ;7708
                                                end
                                                if (((~(P2_P3_r < P2_P3_m)) | (P2_P3_B == 1'b1))) begin
                                                    $display(";A 7710");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))) (bv-comp P2_P3_B  0b1))   0b1)) ;7710
                                                    P2_P3_B = 1'b1; $display(";A 7712");		//(= P2_P3_B    0b1)) ;7712
                                                end
                                                else begin
                                                    $display(";A 7711");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P3_r  P2_P3_m ))) (bv-comp P2_P3_B  0b1))   0b0)) ;7711
                                                    P2_P3_B = 1'b0; $display(";A 7713");		//(= P2_P3_B    0b0)) ;7713
                                                end
                                            end
                                    endcase
                                end
                            1'b0 :
                                begin
                                    $display(";A 7714");		//(= P2_P3_cf    0b0)) ;7714
                                    if ((~(P2_P3_df == 32'b00000000000000000000000000000111))) begin
                                        $display(";A 7715");		//(= (bv-not (bv-comp P2_P3_df  0b00000000000000000000000000000111))   0b1)) ;7715
                                        if ((P2_P3_df == 32'b00000000000000000000000000000101)) begin
                                            $display(";A 7717");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000101)   0b1)) ;7717
                                            if (((~P2_P3_B) == 1'b1)) begin
                                                $display(";A 7719");		//(= (bv-comp (bv-not P2_P3_B ) 0b1)   0b1)) ;7719
                                                P2_P3_d = 32'sb00000000000000000000000000000011; $display(";A 7721");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7721
                                            end
                                            else begin
                                                $display(";A 7720");		//(= (bv-comp (bv-not P2_P3_B ) 0b1)   0b0)) ;7720
                                            end
                                        end
                                        else begin
                                            $display(";A 7718");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000101)   0b0)) ;7718
                                            if ((P2_P3_df == 32'b00000000000000000000000000000100)) begin
                                                $display(";A 7722");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000100)   0b1)) ;7722
                                                if ((P2_P3_B == 1'b1)) begin
                                                    $display(";A 7724");		//(= (bv-comp P2_P3_B  0b1)   0b1)) ;7724
                                                    P2_P3_d = 32'sb00000000000000000000000000000011; $display(";A 7726");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7726
                                                end
                                                else begin
                                                    $display(";A 7725");		//(= (bv-comp P2_P3_B  0b1)   0b0)) ;7725
                                                end
                                            end
                                            else begin
                                                $display(";A 7723");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000100)   0b0)) ;7723
                                                if ((P2_P3_df == 32'b00000000000000000000000000000011)) begin
                                                    $display(";A 7727");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000011)   0b1)) ;7727
                                                    P2_P3_d = 32'sb00000000000000000000000000000011; $display(";A 7729");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7729
                                                end
                                                else begin
                                                    $display(";A 7728");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000011)   0b0)) ;7728
                                                    if ((P2_P3_df == 32'b00000000000000000000000000000010)) begin
                                                        $display(";A 7730");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000010)   0b1)) ;7730
                                                        P2_P3_d = 32'sb00000000000000000000000000000010; $display(";A 7732");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7732
                                                    end
                                                    else begin
                                                        $display(";A 7731");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000010)   0b0)) ;7731
                                                        if ((P2_P3_df == 32'b00000000000000000000000000000001)) begin
                                                            $display(";A 7733");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000001)   0b1)) ;7733
                                                            P2_P3_d = 32'sb00000000000000000000000000000001; $display(";A 7735");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7735
                                                        end
                                                        else begin
                                                            $display(";A 7734");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000001)   0b0)) ;7734
                                                            if ((P2_P3_df == 32'b00000000000000000000000000000000)) begin
                                                                $display(";A 7736");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000000)   0b1)) ;7736
                                                                P2_P3_d = 32'sb00000000000000000000000000000000; $display(";A 7738");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7738
                                                            end
                                                            else begin
                                                                $display(";A 7737");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000000)   0b0)) ;7737
                                                            end
                                                        end
                                                    end
                                                end
                                            end
                                        end
                                        case (P2_P3_ff)
                                            4'b0000 :
                                                begin
                                                    $display(";A 7739");		//(= P2_P3_ff    0b0000)) ;7739
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7740");		//(= P2_P3_mf    0b00)) ;7740
                                                                P2_P3_m = P2_P3_tail; $display(";A 7741");		//(= P2_P3_m    P2_P3_tail )) ;7741
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7742");		//(= P2_P3_mf    0b01)) ;7742
                                                                P2_P3_m = P2_P3_datai; $display(";A 7743");		//(= P2_P3_m    P2_P3_datai )) ;7743
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7744");		//(= P2_P3_addr    P2_P3_tail )) ;7744
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7745");		//(= P2_P3_rd    0b1)) ;7745
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7746");		//(= P2_P3_mf    0b10)) ;7746
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7747");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7747
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7748");		//(= P2_P3_rd    0b1)) ;7748
                                                                P2_P3_m = P2_P3_datai; $display(";A 7749");		//(= P2_P3_m    P2_P3_datai )) ;7749
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7750");		//(= P2_P3_mf    0b11)) ;7750
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7751");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7751
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7752");		//(= P2_P3_rd    0b1)) ;7752
                                                                P2_P3_m = P2_P3_datai; $display(";A 7753");		//(= P2_P3_m    P2_P3_datai )) ;7753
                                                            end
                                                    endcase
                                                    P2_P3_t = 32'sb00000000000000000000000000000000; $display(";A 7754");		//(= P2_P3_t    0b00000000000000000000000000000000)) ;7754
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7755");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7755
                                                                P2_P3_reg0 = (P2_P3_t - P2_P3_m); $display(";A 7756");		//(= P2_P3_reg0    (bv-sub P2_P3_t  P2_P3_m ))) ;7756
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7757");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7757
                                                                P2_P3_reg1 = (P2_P3_t - P2_P3_m); $display(";A 7758");		//(= P2_P3_reg1    (bv-sub P2_P3_t  P2_P3_m ))) ;7758
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7759");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7759
                                                                P2_P3_reg2 = (P2_P3_t - P2_P3_m); $display(";A 7760");		//(= P2_P3_reg2    (bv-sub P2_P3_t  P2_P3_m ))) ;7760
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7761");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7761
                                                                P2_P3_reg3 = (P2_P3_t - P2_P3_m); $display(";A 7762");		//(= P2_P3_reg3    (bv-sub P2_P3_t  P2_P3_m ))) ;7762
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7763");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7763
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0001 :
                                                begin
                                                    $display(";A 7764");		//(= P2_P3_ff    0b0001)) ;7764
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7765");		//(= P2_P3_mf    0b00)) ;7765
                                                                P2_P3_m = P2_P3_tail; $display(";A 7766");		//(= P2_P3_m    P2_P3_tail )) ;7766
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7767");		//(= P2_P3_mf    0b01)) ;7767
                                                                P2_P3_m = P2_P3_datai; $display(";A 7768");		//(= P2_P3_m    P2_P3_datai )) ;7768
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7769");		//(= P2_P3_addr    P2_P3_tail )) ;7769
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7770");		//(= P2_P3_rd    0b1)) ;7770
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7771");		//(= P2_P3_mf    0b10)) ;7771
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7772");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7772
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7773");		//(= P2_P3_rd    0b1)) ;7773
                                                                P2_P3_m = P2_P3_datai; $display(";A 7774");		//(= P2_P3_m    P2_P3_datai )) ;7774
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7775");		//(= P2_P3_mf    0b11)) ;7775
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7776");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7776
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7777");		//(= P2_P3_rd    0b1)) ;7777
                                                                P2_P3_m = P2_P3_datai; $display(";A 7778");		//(= P2_P3_m    P2_P3_datai )) ;7778
                                                            end
                                                    endcase
                                                    P2_P3_reg2 = P2_P3_reg3; $display(";A 7779");		//(= P2_P3_reg2    P2_P3_reg3 )) ;7779
                                                    P2_P3_reg3 = P2_P3_m; $display(";A 7780");		//(= P2_P3_reg3    P2_P3_m )) ;7780
                                                end
                                            4'b0010 :
                                                begin
                                                    $display(";A 7781");		//(= P2_P3_ff    0b0010)) ;7781
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7782");		//(= P2_P3_mf    0b00)) ;7782
                                                                P2_P3_m = P2_P3_tail; $display(";A 7783");		//(= P2_P3_m    P2_P3_tail )) ;7783
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7784");		//(= P2_P3_mf    0b01)) ;7784
                                                                P2_P3_m = P2_P3_datai; $display(";A 7785");		//(= P2_P3_m    P2_P3_datai )) ;7785
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7786");		//(= P2_P3_addr    P2_P3_tail )) ;7786
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7787");		//(= P2_P3_rd    0b1)) ;7787
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7788");		//(= P2_P3_mf    0b10)) ;7788
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7789");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7789
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7790");		//(= P2_P3_rd    0b1)) ;7790
                                                                P2_P3_m = P2_P3_datai; $display(";A 7791");		//(= P2_P3_m    P2_P3_datai )) ;7791
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7792");		//(= P2_P3_mf    0b11)) ;7792
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7793");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7793
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7794");		//(= P2_P3_rd    0b1)) ;7794
                                                                P2_P3_m = P2_P3_datai; $display(";A 7795");		//(= P2_P3_m    P2_P3_datai )) ;7795
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7796");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7796
                                                                P2_P3_reg0 = P2_P3_m; $display(";A 7797");		//(= P2_P3_reg0    P2_P3_m )) ;7797
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7798");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7798
                                                                P2_P3_reg1 = P2_P3_m; $display(";A 7799");		//(= P2_P3_reg1    P2_P3_m )) ;7799
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7800");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7800
                                                                P2_P3_reg2 = P2_P3_m; $display(";A 7801");		//(= P2_P3_reg2    P2_P3_m )) ;7801
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7802");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7802
                                                                P2_P3_reg3 = P2_P3_m; $display(";A 7803");		//(= P2_P3_reg3    P2_P3_m )) ;7803
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7804");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7804
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0011 :
                                                begin
                                                    $display(";A 7805");		//(= P2_P3_ff    0b0011)) ;7805
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7806");		//(= P2_P3_mf    0b00)) ;7806
                                                                P2_P3_m = P2_P3_tail; $display(";A 7807");		//(= P2_P3_m    P2_P3_tail )) ;7807
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7808");		//(= P2_P3_mf    0b01)) ;7808
                                                                P2_P3_m = P2_P3_datai; $display(";A 7809");		//(= P2_P3_m    P2_P3_datai )) ;7809
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7810");		//(= P2_P3_addr    P2_P3_tail )) ;7810
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7811");		//(= P2_P3_rd    0b1)) ;7811
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7812");		//(= P2_P3_mf    0b10)) ;7812
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7813");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7813
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7814");		//(= P2_P3_rd    0b1)) ;7814
                                                                P2_P3_m = P2_P3_datai; $display(";A 7815");		//(= P2_P3_m    P2_P3_datai )) ;7815
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7816");		//(= P2_P3_mf    0b11)) ;7816
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7817");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7817
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7818");		//(= P2_P3_rd    0b1)) ;7818
                                                                P2_P3_m = P2_P3_datai; $display(";A 7819");		//(= P2_P3_m    P2_P3_datai )) ;7819
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7820");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7820
                                                                P2_P3_reg0 = P2_P3_m; $display(";A 7821");		//(= P2_P3_reg0    P2_P3_m )) ;7821
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7822");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7822
                                                                P2_P3_reg1 = P2_P3_m; $display(";A 7823");		//(= P2_P3_reg1    P2_P3_m )) ;7823
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7824");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7824
                                                                P2_P3_reg2 = P2_P3_m; $display(";A 7825");		//(= P2_P3_reg2    P2_P3_m )) ;7825
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7826");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7826
                                                                P2_P3_reg3 = P2_P3_m; $display(";A 7827");		//(= P2_P3_reg3    P2_P3_m )) ;7827
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7828");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7828
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0100 :
                                                begin
                                                    $display(";A 7829");		//(= P2_P3_ff    0b0100)) ;7829
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7830");		//(= P2_P3_mf    0b00)) ;7830
                                                                P2_P3_m = P2_P3_tail; $display(";A 7831");		//(= P2_P3_m    P2_P3_tail )) ;7831
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7832");		//(= P2_P3_mf    0b01)) ;7832
                                                                P2_P3_m = P2_P3_datai; $display(";A 7833");		//(= P2_P3_m    P2_P3_datai )) ;7833
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7834");		//(= P2_P3_addr    P2_P3_tail )) ;7834
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7835");		//(= P2_P3_rd    0b1)) ;7835
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7836");		//(= P2_P3_mf    0b10)) ;7836
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7837");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7837
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7838");		//(= P2_P3_rd    0b1)) ;7838
                                                                P2_P3_m = P2_P3_datai; $display(";A 7839");		//(= P2_P3_m    P2_P3_datai )) ;7839
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7840");		//(= P2_P3_mf    0b11)) ;7840
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7841");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7841
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7842");		//(= P2_P3_rd    0b1)) ;7842
                                                                P2_P3_m = P2_P3_datai; $display(";A 7843");		//(= P2_P3_m    P2_P3_datai )) ;7843
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7844");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7844
                                                                P2_P3_reg0 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7845");		//(= P2_P3_reg0    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7845
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7846");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7846
                                                                P2_P3_reg1 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7847");		//(= P2_P3_reg1    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7847
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7848");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7848
                                                                P2_P3_reg2 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7849");		//(= P2_P3_reg2    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7849
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7850");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7850
                                                                P2_P3_reg3 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7851");		//(= P2_P3_reg3    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7851
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7852");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7852
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0101 :
                                                begin
                                                    $display(";A 7853");		//(= P2_P3_ff    0b0101)) ;7853
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7854");		//(= P2_P3_mf    0b00)) ;7854
                                                                P2_P3_m = P2_P3_tail; $display(";A 7855");		//(= P2_P3_m    P2_P3_tail )) ;7855
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7856");		//(= P2_P3_mf    0b01)) ;7856
                                                                P2_P3_m = P2_P3_datai; $display(";A 7857");		//(= P2_P3_m    P2_P3_datai )) ;7857
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7858");		//(= P2_P3_addr    P2_P3_tail )) ;7858
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7859");		//(= P2_P3_rd    0b1)) ;7859
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7860");		//(= P2_P3_mf    0b10)) ;7860
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7861");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7861
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7862");		//(= P2_P3_rd    0b1)) ;7862
                                                                P2_P3_m = P2_P3_datai; $display(";A 7863");		//(= P2_P3_m    P2_P3_datai )) ;7863
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7864");		//(= P2_P3_mf    0b11)) ;7864
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7865");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7865
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7866");		//(= P2_P3_rd    0b1)) ;7866
                                                                P2_P3_m = P2_P3_datai; $display(";A 7867");		//(= P2_P3_m    P2_P3_datai )) ;7867
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7868");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7868
                                                                P2_P3_reg0 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7869");		//(= P2_P3_reg0    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7869
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7870");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7870
                                                                P2_P3_reg1 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7871");		//(= P2_P3_reg1    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7871
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7872");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7872
                                                                P2_P3_reg2 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7873");		//(= P2_P3_reg2    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7873
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7874");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7874
                                                                P2_P3_reg3 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7875");		//(= P2_P3_reg3    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7875
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7876");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7876
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0110 :
                                                begin
                                                    $display(";A 7877");		//(= P2_P3_ff    0b0110)) ;7877
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7878");		//(= P2_P3_mf    0b00)) ;7878
                                                                P2_P3_m = P2_P3_tail; $display(";A 7879");		//(= P2_P3_m    P2_P3_tail )) ;7879
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7880");		//(= P2_P3_mf    0b01)) ;7880
                                                                P2_P3_m = P2_P3_datai; $display(";A 7881");		//(= P2_P3_m    P2_P3_datai )) ;7881
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7882");		//(= P2_P3_addr    P2_P3_tail )) ;7882
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7883");		//(= P2_P3_rd    0b1)) ;7883
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7884");		//(= P2_P3_mf    0b10)) ;7884
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7885");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7885
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7886");		//(= P2_P3_rd    0b1)) ;7886
                                                                P2_P3_m = P2_P3_datai; $display(";A 7887");		//(= P2_P3_m    P2_P3_datai )) ;7887
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7888");		//(= P2_P3_mf    0b11)) ;7888
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7889");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7889
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7890");		//(= P2_P3_rd    0b1)) ;7890
                                                                P2_P3_m = P2_P3_datai; $display(";A 7891");		//(= P2_P3_m    P2_P3_datai )) ;7891
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7892");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7892
                                                                P2_P3_reg0 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7893");		//(= P2_P3_reg0    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7893
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7894");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7894
                                                                P2_P3_reg1 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7895");		//(= P2_P3_reg1    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7895
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7896");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7896
                                                                P2_P3_reg2 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7897");		//(= P2_P3_reg2    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7897
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7898");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7898
                                                                P2_P3_reg3 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7899");		//(= P2_P3_reg3    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7899
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7900");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7900
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0111 :
                                                begin
                                                    $display(";A 7901");		//(= P2_P3_ff    0b0111)) ;7901
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7902");		//(= P2_P3_mf    0b00)) ;7902
                                                                P2_P3_m = P2_P3_tail; $display(";A 7903");		//(= P2_P3_m    P2_P3_tail )) ;7903
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7904");		//(= P2_P3_mf    0b01)) ;7904
                                                                P2_P3_m = P2_P3_datai; $display(";A 7905");		//(= P2_P3_m    P2_P3_datai )) ;7905
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7906");		//(= P2_P3_addr    P2_P3_tail )) ;7906
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7907");		//(= P2_P3_rd    0b1)) ;7907
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7908");		//(= P2_P3_mf    0b10)) ;7908
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7909");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7909
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7910");		//(= P2_P3_rd    0b1)) ;7910
                                                                P2_P3_m = P2_P3_datai; $display(";A 7911");		//(= P2_P3_m    P2_P3_datai )) ;7911
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7912");		//(= P2_P3_mf    0b11)) ;7912
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7913");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7913
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7914");		//(= P2_P3_rd    0b1)) ;7914
                                                                P2_P3_m = P2_P3_datai; $display(";A 7915");		//(= P2_P3_m    P2_P3_datai )) ;7915
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7916");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7916
                                                                P2_P3_reg0 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7917");		//(= P2_P3_reg0    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7917
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7918");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7918
                                                                P2_P3_reg1 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7919");		//(= P2_P3_reg1    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7919
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7920");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7920
                                                                P2_P3_reg2 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7921");		//(= P2_P3_reg2    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7921
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7922");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7922
                                                                P2_P3_reg3 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7923");		//(= P2_P3_reg3    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7923
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7924");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7924
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1000 :
                                                begin
                                                    $display(";A 7925");		//(= P2_P3_ff    0b1000)) ;7925
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7926");		//(= P2_P3_mf    0b00)) ;7926
                                                                P2_P3_m = P2_P3_tail; $display(";A 7927");		//(= P2_P3_m    P2_P3_tail )) ;7927
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7928");		//(= P2_P3_mf    0b01)) ;7928
                                                                P2_P3_m = P2_P3_datai; $display(";A 7929");		//(= P2_P3_m    P2_P3_datai )) ;7929
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7930");		//(= P2_P3_addr    P2_P3_tail )) ;7930
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7931");		//(= P2_P3_rd    0b1)) ;7931
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7932");		//(= P2_P3_mf    0b10)) ;7932
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7933");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7933
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7934");		//(= P2_P3_rd    0b1)) ;7934
                                                                P2_P3_m = P2_P3_datai; $display(";A 7935");		//(= P2_P3_m    P2_P3_datai )) ;7935
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7936");		//(= P2_P3_mf    0b11)) ;7936
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7937");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7937
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7938");		//(= P2_P3_rd    0b1)) ;7938
                                                                P2_P3_m = P2_P3_datai; $display(";A 7939");		//(= P2_P3_m    P2_P3_datai )) ;7939
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7940");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7940
                                                                P2_P3_reg0 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7941");		//(= P2_P3_reg0    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7941
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7942");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7942
                                                                P2_P3_reg1 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7943");		//(= P2_P3_reg1    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7943
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7944");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7944
                                                                P2_P3_reg2 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7945");		//(= P2_P3_reg2    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7945
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7946");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7946
                                                                P2_P3_reg3 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7947");		//(= P2_P3_reg3    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7947
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7948");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7948
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1001 :
                                                begin
                                                    $display(";A 7949");		//(= P2_P3_ff    0b1001)) ;7949
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7950");		//(= P2_P3_mf    0b00)) ;7950
                                                                P2_P3_m = P2_P3_tail; $display(";A 7951");		//(= P2_P3_m    P2_P3_tail )) ;7951
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7952");		//(= P2_P3_mf    0b01)) ;7952
                                                                P2_P3_m = P2_P3_datai; $display(";A 7953");		//(= P2_P3_m    P2_P3_datai )) ;7953
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7954");		//(= P2_P3_addr    P2_P3_tail )) ;7954
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7955");		//(= P2_P3_rd    0b1)) ;7955
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7956");		//(= P2_P3_mf    0b10)) ;7956
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7957");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7957
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7958");		//(= P2_P3_rd    0b1)) ;7958
                                                                P2_P3_m = P2_P3_datai; $display(";A 7959");		//(= P2_P3_m    P2_P3_datai )) ;7959
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7960");		//(= P2_P3_mf    0b11)) ;7960
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7961");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7961
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7962");		//(= P2_P3_rd    0b1)) ;7962
                                                                P2_P3_m = P2_P3_datai; $display(";A 7963");		//(= P2_P3_m    P2_P3_datai )) ;7963
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7964");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7964
                                                                P2_P3_reg0 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7965");		//(= P2_P3_reg0    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7965
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7966");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7966
                                                                P2_P3_reg1 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7967");		//(= P2_P3_reg1    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7967
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7968");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7968
                                                                P2_P3_reg2 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7969");		//(= P2_P3_reg2    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7969
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7970");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7970
                                                                P2_P3_reg3 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7971");		//(= P2_P3_reg3    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7971
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7972");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7972
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1010 :
                                                begin
                                                    $display(";A 7973");		//(= P2_P3_ff    0b1010)) ;7973
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7974");		//(= P2_P3_mf    0b00)) ;7974
                                                                P2_P3_m = P2_P3_tail; $display(";A 7975");		//(= P2_P3_m    P2_P3_tail )) ;7975
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 7976");		//(= P2_P3_mf    0b01)) ;7976
                                                                P2_P3_m = P2_P3_datai; $display(";A 7977");		//(= P2_P3_m    P2_P3_datai )) ;7977
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 7978");		//(= P2_P3_addr    P2_P3_tail )) ;7978
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7979");		//(= P2_P3_rd    0b1)) ;7979
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 7980");		//(= P2_P3_mf    0b10)) ;7980
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 7981");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;7981
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7982");		//(= P2_P3_rd    0b1)) ;7982
                                                                P2_P3_m = P2_P3_datai; $display(";A 7983");		//(= P2_P3_m    P2_P3_datai )) ;7983
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 7984");		//(= P2_P3_mf    0b11)) ;7984
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 7985");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;7985
                                                                P2_P3_rd <= #1 1'b1; $display(";A 7986");		//(= P2_P3_rd    0b1)) ;7986
                                                                P2_P3_m = P2_P3_datai; $display(";A 7987");		//(= P2_P3_m    P2_P3_datai )) ;7987
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 7988");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;7988
                                                                P2_P3_reg0 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7989");		//(= P2_P3_reg0    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7989
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 7990");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;7990
                                                                P2_P3_reg1 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7991");		//(= P2_P3_reg1    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7991
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 7992");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;7992
                                                                P2_P3_reg2 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7993");		//(= P2_P3_reg2    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7993
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 7994");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;7994
                                                                P2_P3_reg3 = ((P2_P3_r + P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 7995");		//(= P2_P3_reg3    (bv-smod (bv-add P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;7995
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 7996");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;7996
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1011 :
                                                begin
                                                    $display(";A 7997");		//(= P2_P3_ff    0b1011)) ;7997
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 7998");		//(= P2_P3_mf    0b00)) ;7998
                                                                P2_P3_m = P2_P3_tail; $display(";A 7999");		//(= P2_P3_m    P2_P3_tail )) ;7999
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8000");		//(= P2_P3_mf    0b01)) ;8000
                                                                P2_P3_m = P2_P3_datai; $display(";A 8001");		//(= P2_P3_m    P2_P3_datai )) ;8001
                                                                P2_P3_addr <= #1 P2_P3_tail; $display(";A 8002");		//(= P2_P3_addr    P2_P3_tail )) ;8002
                                                                P2_P3_rd <= #1 1'b1; $display(";A 8003");		//(= P2_P3_rd    0b1)) ;8003
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8004");		//(= P2_P3_mf    0b10)) ;8004
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg1) % 32'b00000000000100000000000000000000); $display(";A 8005");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg1 ) 0b00000000000100000000000000000000))) ;8005
                                                                P2_P3_rd <= #1 1'b1; $display(";A 8006");		//(= P2_P3_rd    0b1)) ;8006
                                                                P2_P3_m = P2_P3_datai; $display(";A 8007");		//(= P2_P3_m    P2_P3_datai )) ;8007
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8008");		//(= P2_P3_mf    0b11)) ;8008
                                                                P2_P3_addr <= #1 ((P2_P3_tail + P2_P3_reg2) % 32'b00000000000100000000000000000000); $display(";A 8009");		//(= P2_P3_addr    (bv-smod (bv-add P2_P3_tail  P2_P3_reg2 ) 0b00000000000100000000000000000000))) ;8009
                                                                P2_P3_rd <= #1 1'b1; $display(";A 8010");		//(= P2_P3_rd    0b1)) ;8010
                                                                P2_P3_m = P2_P3_datai; $display(";A 8011");		//(= P2_P3_m    P2_P3_datai )) ;8011
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8012");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;8012
                                                                P2_P3_reg0 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 8013");		//(= P2_P3_reg0    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;8013
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8014");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;8014
                                                                P2_P3_reg1 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 8015");		//(= P2_P3_reg1    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;8015
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8016");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;8016
                                                                P2_P3_reg2 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 8017");		//(= P2_P3_reg2    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;8017
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8018");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;8018
                                                                P2_P3_reg3 = ((P2_P3_r - P2_P3_m) % 32'b00000000000000000000000000000000); $display(";A 8019");		//(= P2_P3_reg3    (bv-smod (bv-sub P2_P3_r  P2_P3_m ) 0b00000000000000000000000000000000))) ;8019
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8020");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;8020
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1100 :
                                                begin
                                                    $display(";A 8021");		//(= P2_P3_ff    0b1100)) ;8021
                                                    case (P2_P3_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8022");		//(= P2_P3_mf    0b00)) ;8022
                                                                P2_P3_t = (P2_P3_r / 32'sb00000000000000000000000000000010); $display(";A 8023");		//(= P2_P3_t    (bv-sdiv P2_P3_r  0b00000000000000000000000000000010))) ;8023
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8024");		//(= P2_P3_mf    0b01)) ;8024
                                                                P2_P3_t = (P2_P3_r / 32'sb00000000000000000000000000000010); $display(";A 8025");		//(= P2_P3_t    (bv-sdiv P2_P3_r  0b00000000000000000000000000000010))) ;8025
                                                                if ((P2_P3_B == 1'b1)) begin
                                                                    $display(";A 8026");		//(= (bv-comp P2_P3_B  0b1)   0b1)) ;8026
                                                                    P2_P3_t = (P2_P3_t % 32'b00100000000000000000000000000000); $display(";A 8028");		//(= P2_P3_t    (bv-smod P2_P3_t  0b00100000000000000000000000000000))) ;8028
                                                                end
                                                                else begin
                                                                    $display(";A 8027");		//(= (bv-comp P2_P3_B  0b1)   0b0)) ;8027
                                                                end
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8029");		//(= P2_P3_mf    0b10)) ;8029
                                                                P2_P3_t = ((P2_P3_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 8030");		//(= P2_P3_t    (bv-mul (bv-smod P2_P3_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;8030
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8031");		//(= P2_P3_mf    0b11)) ;8031
                                                                P2_P3_t = ((P2_P3_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 8032");		//(= P2_P3_t    (bv-mul (bv-smod P2_P3_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;8032
                                                                if ((P2_P3_t > 32'b11111111111111111111111111111111)) begin
                                                                    $display(";A 8033");		//(= (bool-to-bv (bv-gt P2_P3_t  0b11111111111111111111111111111111))   0b1)) ;8033
                                                                    P2_P3_B = 1'b1; $display(";A 8035");		//(= P2_P3_B    0b1)) ;8035
                                                                end
                                                                else begin
                                                                    $display(";A 8034");		//(= (bool-to-bv (bv-gt P2_P3_t  0b11111111111111111111111111111111))   0b0)) ;8034
                                                                    P2_P3_B = 1'b0; $display(";A 8036");		//(= P2_P3_B    0b0)) ;8036
                                                                end
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8037");		//(= (and (/= P2_P3_mf  0b00) (/= P2_P3_mf  0b01) (/= P2_P3_mf  0b10) (/= P2_P3_mf  0b11))   true)) ;8037
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                    case (P2_P3_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8038");		//(= P2_P3_d    0b00000000000000000000000000000000)) ;8038
                                                                P2_P3_reg0 = P2_P3_t; $display(";A 8039");		//(= P2_P3_reg0    P2_P3_t )) ;8039
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8040");		//(= P2_P3_d    0b00000000000000000000000000000001)) ;8040
                                                                P2_P3_reg1 = P2_P3_t; $display(";A 8041");		//(= P2_P3_reg1    P2_P3_t )) ;8041
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8042");		//(= P2_P3_d    0b00000000000000000000000000000010)) ;8042
                                                                P2_P3_reg2 = P2_P3_t; $display(";A 8043");		//(= P2_P3_reg2    P2_P3_t )) ;8043
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8044");		//(= P2_P3_d    0b00000000000000000000000000000011)) ;8044
                                                                P2_P3_reg3 = P2_P3_t; $display(";A 8045");		//(= P2_P3_reg3    P2_P3_t )) ;8045
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8046");		//(= (and (/= P2_P3_d  0b00000000000000000000000000000000) (/= P2_P3_d  0b00000000000000000000000000000001) (/= P2_P3_d  0b00000000000000000000000000000010) (/= P2_P3_d  0b00000000000000000000000000000011))   true)) ;8046
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1101 :
                                                begin
                                                    $display(";A 8047");		//(= P2_P3_ff    0b1101)) ;8047
                                                    begin
                                                    end
                                                end
                                            4'b1110 :
                                                begin
                                                    $display(";A 8048");		//(= P2_P3_ff    0b1110)) ;8048
                                                    begin
                                                    end
                                                end
                                            4'b1111 :
                                                begin
                                                    $display(";A 8049");		//(= P2_P3_ff    0b1111)) ;8049
                                                    begin
                                                    end
                                                end
                                        endcase
                                    end
                                    else begin
                                        $display(";A 7716");		//(= (bv-not (bv-comp P2_P3_df  0b00000000000000000000000000000111))   0b0)) ;7716
                                        if ((P2_P3_df == 32'b00000000000000000000000000000111)) begin
                                            $display(";A 8050");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000111)   0b1)) ;8050
                                            case (P2_P3_mf)
                                                2'b00 :
                                                    begin
                                                        $display(";A 8052");		//(= P2_P3_mf    0b00)) ;8052
                                                        P2_P3_m = P2_P3_tail; $display(";A 8053");		//(= P2_P3_m    P2_P3_tail )) ;8053
                                                    end
                                                2'b01 :
                                                    begin
                                                        $display(";A 8054");		//(= P2_P3_mf    0b01)) ;8054
                                                        P2_P3_m = P2_P3_tail; $display(";A 8055");		//(= P2_P3_m    P2_P3_tail )) ;8055
                                                    end
                                                2'b10 :
                                                    begin
                                                        $display(";A 8056");		//(= P2_P3_mf    0b10)) ;8056
                                                        P2_P3_m = ((P2_P3_reg1 % 32'b00000000000100000000000000000000) + (P2_P3_tail % 32'b00000000000100000000000000000000)); $display(";A 8057");		//(= P2_P3_m    (bv-add (bv-smod P2_P3_reg1  0b00000000000100000000000000000000) (bv-smod P2_P3_tail  0b00000000000100000000000000000000)))) ;8057
                                                    end
                                                2'b11 :
                                                    begin
                                                        $display(";A 8058");		//(= P2_P3_mf    0b11)) ;8058
                                                        P2_P3_m = ((P2_P3_reg2 % 32'b00000000000100000000000000000000) + (P2_P3_tail % 32'b00000000000100000000000000000000)); $display(";A 8059");		//(= P2_P3_m    (bv-add (bv-smod P2_P3_reg2  0b00000000000100000000000000000000) (bv-smod P2_P3_tail  0b00000000000100000000000000000000)))) ;8059
                                                    end
                                            endcase
                                            P2_P3_addr <= #1 ((P2_P3_m % 32'sb00000000000000000000000000000010) * 32'sb00000000000000000000000000010100); $display(";A 8060");		//(= P2_P3_addr    (bv-mul (bv-smod P2_P3_m  0b00000000000000000000000000000010) 0b00000000000000000000000000010100))) ;8060
                                            P2_P3_wr <= #1 1'b1; $display(";A 8061");		//(= P2_P3_wr    0b1)) ;8061
                                            P2_P3_datao <= #1 P2_P3_r; $display(";A 8062");		//(= P2_P3_datao    P2_P3_r )) ;8062
                                        end
                                        else begin
                                            $display(";A 8051");		//(= (bv-comp P2_P3_df  0b00000000000000000000000000000111)   0b0)) ;8051
                                        end
                                    end
                                end
                        endcase
                        P2_P3_state = 1'sb0; $display(";A 8063");		//(= P2_P3_state    0b0)) ;8063
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:12357
    always @(posedge P2_P4_reset or posedge P2_P4_clock) begin
        if ((P2_P4_reset == 1'b1)) begin
            P2_P4_MAR = 20'sb00000000000000000000; $display(";A 8066");		//(= P2_P4_MAR    0b00000000000000000000)) ;8066
            P2_P4_MBR = 32'sb00000000000000000000000000000000; $display(";A 8067");		//(= P2_P4_MBR    0b00000000000000000000000000000000)) ;8067
            P2_P4_IR = 32'sb00000000000000000000000000000000; $display(";A 8068");		//(= P2_P4_IR    0b00000000000000000000000000000000)) ;8068
            P2_P4_d = 32'sb00000000000000000000000000000000; $display(";A 8069");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8069
            P2_P4_r = 32'sb00000000000000000000000000000000; $display(";A 8070");		//(= P2_P4_r    0b00000000000000000000000000000000)) ;8070
            P2_P4_m = 32'sb00000000000000000000000000000000; $display(";A 8071");		//(= P2_P4_m    0b00000000000000000000000000000000)) ;8071
            P2_P4_s = 2'sb00; $display(";A 8072");		//(= P2_P4_s    0b00)) ;8072
            P2_P4_temp = 32'sb00000000000000000000000000000000; $display(";A 8073");		//(= P2_P4_temp    0b00000000000000000000000000000000)) ;8073
            P2_P4_mf = 2'sb00; $display(";A 8074");		//(= P2_P4_mf    0b00)) ;8074
            P2_P4_df = 3'sb000; $display(";A 8075");		//(= P2_P4_df    0b000)) ;8075
            P2_P4_ff = 4'sb0000; $display(";A 8076");		//(= P2_P4_ff    0b0000)) ;8076
            P2_P4_cf = 1'sb0; $display(";A 8077");		//(= P2_P4_cf    0b0)) ;8077
            P2_P4_tail = 20'sb00000000000000000000; $display(";A 8078");		//(= P2_P4_tail    0b00000000000000000000)) ;8078
            P2_P4_B = 1'b0; $display(";A 8079");		//(= P2_P4_B    0b0)) ;8079
            P2_P4_reg0 = 32'sb00000000000000000000000000000000; $display(";A 8080");		//(= P2_P4_reg0    0b00000000000000000000000000000000)) ;8080
            P2_P4_reg1 = 32'sb00000000000000000000000000000000; $display(";A 8081");		//(= P2_P4_reg1    0b00000000000000000000000000000000)) ;8081
            P2_P4_reg2 = 32'sb00000000000000000000000000000000; $display(";A 8082");		//(= P2_P4_reg2    0b00000000000000000000000000000000)) ;8082
            P2_P4_reg3 = 32'sb00000000000000000000000000000000; $display(";A 8083");		//(= P2_P4_reg3    0b00000000000000000000000000000000)) ;8083
            P2_P4_addr <= #1 20'sb00000000000000000000; $display(";A 8084");		//(= P2_P4_addr    0b00000000000000000000)) ;8084
            P2_P4_rd <= #1 1'b0; $display(";A 8085");		//(= P2_P4_rd    0b0)) ;8085
            P2_P4_wr <= #1 1'b0; $display(";A 8086");		//(= P2_P4_wr    0b0)) ;8086
            P2_P4_datao <= #1 32'sb00000000000000000000000000000000; $display(";A 8087");		//(= P2_P4_datao    0b00000000000000000000000000000000)) ;8087
            P2_P4_state = 1'sb0; $display(";A 8088");		//(= P2_P4_state    0b0)) ;8088
        end
        else begin
            P2_P4_rd <= #1 1'b0; $display(";A 8089");		//(= P2_P4_rd    0b0)) ;8089
            P2_P4_wr <= #1 1'b0; $display(";A 8090");		//(= P2_P4_wr    0b0)) ;8090
            case (P2_P4_state)
                1'b0 :
                    begin
                        $display(";A 8091");		//(= P2_P4_state    0b0)) ;8091
                        P2_P4_MAR = (P2_P4_reg3 % 32'b00000000000100000000000000000000); $display(";A 8092");		//(= P2_P4_MAR    (bv-smod P2_P4_reg3  0b00000000000100000000000000000000))) ;8092
                        P2_P4_addr <= #1 P2_P4_MAR; $display(";A 8093");		//(= P2_P4_addr    P2_P4_MAR )) ;8093
                        P2_P4_rd <= #1 1'b1; $display(";A 8094");		//(= P2_P4_rd    0b1)) ;8094
                        P2_P4_MBR = P2_P4_datai; $display(";A 8095");		//(= P2_P4_MBR    P2_P4_datai )) ;8095
                        P2_P4_IR = P2_P4_MBR; $display(";A 8096");		//(= P2_P4_IR    P2_P4_MBR )) ;8096
                        P2_P4_state = 1'sb1; $display(";A 8097");		//(= P2_P4_state    0b1)) ;8097
                    end
                1'b1 :
                    begin
                        $display(";A 8098");		//(= P2_P4_state    0b1)) ;8098
                        if ((P2_P4_IR < 32'sb00000000000000000000000000000000)) begin
                            $display(";A 8099");		//(= (bool-to-bv (bv-slt P2_P4_IR  0b00000000000000000000000000000000))   0b1)) ;8099
                            P2_P4_IR = (-P2_P4_IR); $display(";A 8101");		//(= P2_P4_IR    (bv-neg P2_P4_IR ))) ;8101
                        end
                        else begin
                            $display(";A 8100");		//(= (bool-to-bv (bv-slt P2_P4_IR  0b00000000000000000000000000000000))   0b0)) ;8100
                        end
                        P2_P4_mf = ((P2_P4_IR / 32'b00001000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 8102");		//(= P2_P4_mf    (bv-smod (bv-sdiv P2_P4_IR  0b00001000000000000000000000000000) 0b00000000000000000000000000000100))) ;8102
                        P2_P4_df = ((P2_P4_IR / 32'b00000001000000000000000000000000) % 32'b00000000000000000000000000001000); $display(";A 8103");		//(= P2_P4_df    (bv-smod (bv-sdiv P2_P4_IR  0b00000001000000000000000000000000) 0b00000000000000000000000000001000))) ;8103
                        P2_P4_ff = ((P2_P4_IR / 32'b00000000000010000000000000000000) % 32'b00000000000000000000000000010000); $display(";A 8104");		//(= P2_P4_ff    (bv-smod (bv-sdiv P2_P4_IR  0b00000000000010000000000000000000) 0b00000000000000000000000000010000))) ;8104
                        P2_P4_cf = ((P2_P4_IR / 32'b00000000100000000000000000000000) % 32'b00000000000000000000000000000010); $display(";A 8105");		//(= P2_P4_cf    (bv-smod (bv-sdiv P2_P4_IR  0b00000000100000000000000000000000) 0b00000000000000000000000000000010))) ;8105
                        P2_P4_tail = (P2_P4_IR % 32'b00000000000100000000000000000000); $display(";A 8106");		//(= P2_P4_tail    (bv-smod P2_P4_IR  0b00000000000100000000000000000000))) ;8106
                        P2_P4_reg3 = ((P2_P4_reg3 % 32'b00100000000000000000000000000000) + 32'b00000000000000000000000000001000); $display(";A 8107");		//(= P2_P4_reg3    (bv-add (bv-smod P2_P4_reg3  0b00100000000000000000000000000000) 0b00000000000000000000000000001000))) ;8107
                        P2_P4_s = ((P2_P4_IR / 32'b00100000000000000000000000000000) % 32'b00000000000000000000000000000100); $display(";A 8108");		//(= P2_P4_s    (bv-smod (bv-sdiv P2_P4_IR  0b00100000000000000000000000000000) 0b00000000000000000000000000000100))) ;8108
                        case (P2_P4_s)
                            2'b00 :
                                begin
                                    $display(";A 8109");		//(= P2_P4_s    0b00)) ;8109
                                    P2_P4_r = P2_P4_reg0; $display(";A 8110");		//(= P2_P4_r    P2_P4_reg0 )) ;8110
                                end
                            2'b01 :
                                begin
                                    $display(";A 8111");		//(= P2_P4_s    0b01)) ;8111
                                    P2_P4_r = P2_P4_reg1; $display(";A 8112");		//(= P2_P4_r    P2_P4_reg1 )) ;8112
                                end
                            2'b10 :
                                begin
                                    $display(";A 8113");		//(= P2_P4_s    0b10)) ;8113
                                    P2_P4_r = P2_P4_reg2; $display(";A 8114");		//(= P2_P4_r    P2_P4_reg2 )) ;8114
                                end
                            2'b11 :
                                begin
                                    $display(";A 8115");		//(= P2_P4_s    0b11)) ;8115
                                    P2_P4_r = P2_P4_reg3; $display(";A 8116");		//(= P2_P4_r    P2_P4_reg3 )) ;8116
                                end
                        endcase
                        case (P2_P4_cf)
                            1'b1 :
                                begin
                                    $display(";A 8117");		//(= P2_P4_cf    0b1)) ;8117
                                    case (P2_P4_mf)
                                        2'b00 :
                                            begin
                                                $display(";A 8118");		//(= P2_P4_mf    0b00)) ;8118
                                                P2_P4_m = P2_P4_tail; $display(";A 8119");		//(= P2_P4_m    P2_P4_tail )) ;8119
                                            end
                                        2'b01 :
                                            begin
                                                $display(";A 8120");		//(= P2_P4_mf    0b01)) ;8120
                                                P2_P4_m = P2_P4_datai; $display(";A 8121");		//(= P2_P4_m    P2_P4_datai )) ;8121
                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8122");		//(= P2_P4_addr    P2_P4_tail )) ;8122
                                                P2_P4_rd <= #1 1'b1; $display(";A 8123");		//(= P2_P4_rd    0b1)) ;8123
                                            end
                                        2'b10 :
                                            begin
                                                $display(";A 8124");		//(= P2_P4_mf    0b10)) ;8124
                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8125");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8125
                                                P2_P4_rd <= #1 1'b1; $display(";A 8126");		//(= P2_P4_rd    0b1)) ;8126
                                                P2_P4_m = P2_P4_datai; $display(";A 8127");		//(= P2_P4_m    P2_P4_datai )) ;8127
                                            end
                                        2'b11 :
                                            begin
                                                $display(";A 8128");		//(= P2_P4_mf    0b11)) ;8128
                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8129");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8129
                                                P2_P4_rd <= #1 1'b1; $display(";A 8130");		//(= P2_P4_rd    0b1)) ;8130
                                                P2_P4_m = P2_P4_datai; $display(";A 8131");		//(= P2_P4_m    P2_P4_datai )) ;8131
                                            end
                                    endcase
                                    case (P2_P4_ff)
                                        4'b0000 :
                                            begin
                                                $display(";A 8132");		//(= P2_P4_ff    0b0000)) ;8132
                                                if ((P2_P4_r < P2_P4_m)) begin
                                                    $display(";A 8133");		//(= (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))   0b1)) ;8133
                                                    P2_P4_B = 1'b1; $display(";A 8135");		//(= P2_P4_B    0b1)) ;8135
                                                end
                                                else begin
                                                    $display(";A 8134");		//(= (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))   0b0)) ;8134
                                                    P2_P4_B = 1'b0; $display(";A 8136");		//(= P2_P4_B    0b0)) ;8136
                                                end
                                            end
                                        4'b0001 :
                                            begin
                                                $display(";A 8137");		//(= P2_P4_ff    0b0001)) ;8137
                                                if ((~(P2_P4_r < P2_P4_m))) begin
                                                    $display(";A 8138");		//(= (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )))   0b1)) ;8138
                                                    P2_P4_B = 1'b1; $display(";A 8140");		//(= P2_P4_B    0b1)) ;8140
                                                end
                                                else begin
                                                    $display(";A 8139");		//(= (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )))   0b0)) ;8139
                                                    P2_P4_B = 1'b0; $display(";A 8141");		//(= P2_P4_B    0b0)) ;8141
                                                end
                                            end
                                        4'b0010 :
                                            begin
                                                $display(";A 8142");		//(= P2_P4_ff    0b0010)) ;8142
                                                if ((P2_P4_r == P2_P4_m)) begin
                                                    $display(";A 8143");		//(= (bv-comp P2_P4_r  P2_P4_m )   0b1)) ;8143
                                                    P2_P4_B = 1'b1; $display(";A 8145");		//(= P2_P4_B    0b1)) ;8145
                                                end
                                                else begin
                                                    $display(";A 8144");		//(= (bv-comp P2_P4_r  P2_P4_m )   0b0)) ;8144
                                                    P2_P4_B = 1'b0; $display(";A 8146");		//(= P2_P4_B    0b0)) ;8146
                                                end
                                            end
                                        4'b0011 :
                                            begin
                                                $display(";A 8147");		//(= P2_P4_ff    0b0011)) ;8147
                                                if ((~(P2_P4_r == P2_P4_m))) begin
                                                    $display(";A 8148");		//(= (bv-not (bv-comp P2_P4_r  P2_P4_m ))   0b1)) ;8148
                                                    P2_P4_B = 1'b1; $display(";A 8150");		//(= P2_P4_B    0b1)) ;8150
                                                end
                                                else begin
                                                    $display(";A 8149");		//(= (bv-not (bv-comp P2_P4_r  P2_P4_m ))   0b0)) ;8149
                                                    P2_P4_B = 1'b0; $display(";A 8151");		//(= P2_P4_B    0b0)) ;8151
                                                end
                                            end
                                        4'b0100 :
                                            begin
                                                $display(";A 8152");		//(= P2_P4_ff    0b0100)) ;8152
                                                if ((~(P2_P4_r > P2_P4_m))) begin
                                                    $display(";A 8153");		//(= (bv-not (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m )))   0b1)) ;8153
                                                    P2_P4_B = 1'b1; $display(";A 8155");		//(= P2_P4_B    0b1)) ;8155
                                                end
                                                else begin
                                                    $display(";A 8154");		//(= (bv-not (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m )))   0b0)) ;8154
                                                    P2_P4_B = 1'b0; $display(";A 8156");		//(= P2_P4_B    0b0)) ;8156
                                                end
                                            end
                                        4'b0101 :
                                            begin
                                                $display(";A 8157");		//(= P2_P4_ff    0b0101)) ;8157
                                                if ((P2_P4_r > P2_P4_m)) begin
                                                    $display(";A 8158");		//(= (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m ))   0b1)) ;8158
                                                    P2_P4_B = 1'b1; $display(";A 8160");		//(= P2_P4_B    0b1)) ;8160
                                                end
                                                else begin
                                                    $display(";A 8159");		//(= (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m ))   0b0)) ;8159
                                                    P2_P4_B = 1'b0; $display(";A 8161");		//(= P2_P4_B    0b0)) ;8161
                                                end
                                            end
                                        4'b0110 :
                                            begin
                                                $display(";A 8162");		//(= P2_P4_ff    0b0110)) ;8162
                                                if ((P2_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 8163");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b1)) ;8163
                                                    P2_P4_r = (P2_P4_r - 32'b00000000000000000000000000000000); $display(";A 8165");		//(= P2_P4_r    (bv-sub P2_P4_r  0b00000000000000000000000000000000))) ;8165
                                                end
                                                else begin
                                                    $display(";A 8164");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b0)) ;8164
                                                end
                                                if ((P2_P4_r < P2_P4_m)) begin
                                                    $display(";A 8166");		//(= (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))   0b1)) ;8166
                                                    P2_P4_B = 1'b1; $display(";A 8168");		//(= P2_P4_B    0b1)) ;8168
                                                end
                                                else begin
                                                    $display(";A 8167");		//(= (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))   0b0)) ;8167
                                                    P2_P4_B = 1'b0; $display(";A 8169");		//(= P2_P4_B    0b0)) ;8169
                                                end
                                            end
                                        4'b0111 :
                                            begin
                                                $display(";A 8170");		//(= P2_P4_ff    0b0111)) ;8170
                                                if ((P2_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 8171");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b1)) ;8171
                                                    P2_P4_r = (P2_P4_r - 32'b00000000000000000000000000000000); $display(";A 8173");		//(= P2_P4_r    (bv-sub P2_P4_r  0b00000000000000000000000000000000))) ;8173
                                                end
                                                else begin
                                                    $display(";A 8172");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b0)) ;8172
                                                end
                                                if ((~(P2_P4_r < P2_P4_m))) begin
                                                    $display(";A 8174");		//(= (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )))   0b1)) ;8174
                                                    P2_P4_B = 1'b1; $display(";A 8176");		//(= P2_P4_B    0b1)) ;8176
                                                end
                                                else begin
                                                    $display(";A 8175");		//(= (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )))   0b0)) ;8175
                                                    P2_P4_B = 1'b0; $display(";A 8177");		//(= P2_P4_B    0b0)) ;8177
                                                end
                                            end
                                        4'b1000 :
                                            begin
                                                $display(";A 8178");		//(= P2_P4_ff    0b1000)) ;8178
                                                if (((P2_P4_r < P2_P4_m) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8179");		//(= (bv-or (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b1)) ;8179
                                                    P2_P4_B = 1'b1; $display(";A 8181");		//(= P2_P4_B    0b1)) ;8181
                                                end
                                                else begin
                                                    $display(";A 8180");		//(= (bv-or (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b0)) ;8180
                                                    P2_P4_B = 1'b0; $display(";A 8182");		//(= P2_P4_B    0b0)) ;8182
                                                end
                                            end
                                        4'b1001 :
                                            begin
                                                $display(";A 8183");		//(= P2_P4_ff    0b1001)) ;8183
                                                if (((~(P2_P4_r < P2_P4_m)) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8184");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))) (bv-comp P2_P4_B  0b1))   0b1)) ;8184
                                                    P2_P4_B = 1'b1; $display(";A 8186");		//(= P2_P4_B    0b1)) ;8186
                                                end
                                                else begin
                                                    $display(";A 8185");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))) (bv-comp P2_P4_B  0b1))   0b0)) ;8185
                                                    P2_P4_B = 1'b0; $display(";A 8187");		//(= P2_P4_B    0b0)) ;8187
                                                end
                                            end
                                        4'b1010 :
                                            begin
                                                $display(";A 8188");		//(= P2_P4_ff    0b1010)) ;8188
                                                if (((P2_P4_r == P2_P4_m) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8189");		//(= (bv-or (bv-comp P2_P4_r  P2_P4_m ) (bv-comp P2_P4_B  0b1))   0b1)) ;8189
                                                    P2_P4_B = 1'b1; $display(";A 8191");		//(= P2_P4_B    0b1)) ;8191
                                                end
                                                else begin
                                                    $display(";A 8190");		//(= (bv-or (bv-comp P2_P4_r  P2_P4_m ) (bv-comp P2_P4_B  0b1))   0b0)) ;8190
                                                    P2_P4_B = 1'b0; $display(";A 8192");		//(= P2_P4_B    0b0)) ;8192
                                                end
                                            end
                                        4'b1011 :
                                            begin
                                                $display(";A 8193");		//(= P2_P4_ff    0b1011)) ;8193
                                                if (((~(P2_P4_r == P2_P4_m)) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8194");		//(= (bv-or (bv-not (bv-comp P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b1)) ;8194
                                                    P2_P4_B = 1'b1; $display(";A 8196");		//(= P2_P4_B    0b1)) ;8196
                                                end
                                                else begin
                                                    $display(";A 8195");		//(= (bv-or (bv-not (bv-comp P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b0)) ;8195
                                                    P2_P4_B = 1'b0; $display(";A 8197");		//(= P2_P4_B    0b0)) ;8197
                                                end
                                            end
                                        4'b1100 :
                                            begin
                                                $display(";A 8198");		//(= P2_P4_ff    0b1100)) ;8198
                                                if (((~(P2_P4_r > P2_P4_m)) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8199");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m ))) (bv-comp P2_P4_B  0b1))   0b1)) ;8199
                                                    P2_P4_B = 1'b1; $display(";A 8201");		//(= P2_P4_B    0b1)) ;8201
                                                end
                                                else begin
                                                    $display(";A 8200");		//(= (bv-or (bv-not (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m ))) (bv-comp P2_P4_B  0b1))   0b0)) ;8200
                                                    P2_P4_B = 1'b0; $display(";A 8202");		//(= P2_P4_B    0b0)) ;8202
                                                end
                                            end
                                        4'b1101 :
                                            begin
                                                $display(";A 8203");		//(= P2_P4_ff    0b1101)) ;8203
                                                if (((P2_P4_r > P2_P4_m) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8204");		//(= (bv-or (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b1)) ;8204
                                                    P2_P4_B = 1'b1; $display(";A 8206");		//(= P2_P4_B    0b1)) ;8206
                                                end
                                                else begin
                                                    $display(";A 8205");		//(= (bv-or (bool-to-bv (bv-sgt P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b0)) ;8205
                                                    P2_P4_B = 1'b0; $display(";A 8207");		//(= P2_P4_B    0b0)) ;8207
                                                end
                                            end
                                        4'b1110 :
                                            begin
                                                $display(";A 8208");		//(= P2_P4_ff    0b1110)) ;8208
                                                if ((P2_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 8209");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b1)) ;8209
                                                    P2_P4_r = (P2_P4_r - 32'b00000000000000000000000000000000); $display(";A 8211");		//(= P2_P4_r    (bv-sub P2_P4_r  0b00000000000000000000000000000000))) ;8211
                                                end
                                                else begin
                                                    $display(";A 8210");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b0)) ;8210
                                                end
                                                if (((P2_P4_r < P2_P4_m) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8212");		//(= (bv-or (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b1)) ;8212
                                                    P2_P4_B = 1'b1; $display(";A 8214");		//(= P2_P4_B    0b1)) ;8214
                                                end
                                                else begin
                                                    $display(";A 8213");		//(= (bv-or (bool-to-bv (bv-slt P2_P4_r  P2_P4_m )) (bv-comp P2_P4_B  0b1))   0b0)) ;8213
                                                    P2_P4_B = 1'b0; $display(";A 8215");		//(= P2_P4_B    0b0)) ;8215
                                                end
                                            end
                                        4'b1111 :
                                            begin
                                                $display(";A 8216");		//(= P2_P4_ff    0b1111)) ;8216
                                                if ((P2_P4_r > 32'b11111111111111111111111111111111)) begin
                                                    $display(";A 8217");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b1)) ;8217
                                                    P2_P4_r = (P2_P4_r - 32'b00000000000000000000000000000000); $display(";A 8219");		//(= P2_P4_r    (bv-sub P2_P4_r  0b00000000000000000000000000000000))) ;8219
                                                end
                                                else begin
                                                    $display(";A 8218");		//(= (bool-to-bv (bv-gt P2_P4_r  0b11111111111111111111111111111111))   0b0)) ;8218
                                                end
                                                if (((~(P2_P4_r < P2_P4_m)) | (P2_P4_B == 1'b1))) begin
                                                    $display(";A 8220");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))) (bv-comp P2_P4_B  0b1))   0b1)) ;8220
                                                    P2_P4_B = 1'b1; $display(";A 8222");		//(= P2_P4_B    0b1)) ;8222
                                                end
                                                else begin
                                                    $display(";A 8221");		//(= (bv-or (bv-not (bool-to-bv (bv-slt P2_P4_r  P2_P4_m ))) (bv-comp P2_P4_B  0b1))   0b0)) ;8221
                                                    P2_P4_B = 1'b0; $display(";A 8223");		//(= P2_P4_B    0b0)) ;8223
                                                end
                                            end
                                    endcase
                                end
                            1'b0 :
                                begin
                                    $display(";A 8224");		//(= P2_P4_cf    0b0)) ;8224
                                    if ((~(P2_P4_df == 32'b00000000000000000000000000000111))) begin
                                        $display(";A 8225");		//(= (bv-not (bv-comp P2_P4_df  0b00000000000000000000000000000111))   0b1)) ;8225
                                        if ((P2_P4_df == 32'b00000000000000000000000000000101)) begin
                                            $display(";A 8227");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000101)   0b1)) ;8227
                                            if (((~P2_P4_B) == 1'b1)) begin
                                                $display(";A 8229");		//(= (bv-comp (bv-not P2_P4_B ) 0b1)   0b1)) ;8229
                                                P2_P4_d = 32'sb00000000000000000000000000000011; $display(";A 8231");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8231
                                            end
                                            else begin
                                                $display(";A 8230");		//(= (bv-comp (bv-not P2_P4_B ) 0b1)   0b0)) ;8230
                                            end
                                        end
                                        else begin
                                            $display(";A 8228");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000101)   0b0)) ;8228
                                            if ((P2_P4_df == 32'b00000000000000000000000000000100)) begin
                                                $display(";A 8232");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000100)   0b1)) ;8232
                                                if ((P2_P4_B == 1'b1)) begin
                                                    $display(";A 8234");		//(= (bv-comp P2_P4_B  0b1)   0b1)) ;8234
                                                    P2_P4_d = 32'sb00000000000000000000000000000011; $display(";A 8236");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8236
                                                end
                                                else begin
                                                    $display(";A 8235");		//(= (bv-comp P2_P4_B  0b1)   0b0)) ;8235
                                                end
                                            end
                                            else begin
                                                $display(";A 8233");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000100)   0b0)) ;8233
                                                if ((P2_P4_df == 32'b00000000000000000000000000000011)) begin
                                                    $display(";A 8237");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000011)   0b1)) ;8237
                                                    P2_P4_d = 32'sb00000000000000000000000000000011; $display(";A 8239");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8239
                                                end
                                                else begin
                                                    $display(";A 8238");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000011)   0b0)) ;8238
                                                    if ((P2_P4_df == 32'b00000000000000000000000000000010)) begin
                                                        $display(";A 8240");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000010)   0b1)) ;8240
                                                        P2_P4_d = 32'sb00000000000000000000000000000010; $display(";A 8242");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8242
                                                    end
                                                    else begin
                                                        $display(";A 8241");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000010)   0b0)) ;8241
                                                        if ((P2_P4_df == 32'b00000000000000000000000000000001)) begin
                                                            $display(";A 8243");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000001)   0b1)) ;8243
                                                            P2_P4_d = 32'sb00000000000000000000000000000001; $display(";A 8245");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8245
                                                        end
                                                        else begin
                                                            $display(";A 8244");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000001)   0b0)) ;8244
                                                            if ((P2_P4_df == 32'b00000000000000000000000000000000)) begin
                                                                $display(";A 8246");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000000)   0b1)) ;8246
                                                                P2_P4_d = 32'sb00000000000000000000000000000000; $display(";A 8248");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8248
                                                            end
                                                            else begin
                                                                $display(";A 8247");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000000)   0b0)) ;8247
                                                            end
                                                        end
                                                    end
                                                end
                                            end
                                        end
                                        case (P2_P4_ff)
                                            4'b0000 :
                                                begin
                                                    $display(";A 8249");		//(= P2_P4_ff    0b0000)) ;8249
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8250");		//(= P2_P4_mf    0b00)) ;8250
                                                                P2_P4_m = P2_P4_tail; $display(";A 8251");		//(= P2_P4_m    P2_P4_tail )) ;8251
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8252");		//(= P2_P4_mf    0b01)) ;8252
                                                                P2_P4_m = P2_P4_datai; $display(";A 8253");		//(= P2_P4_m    P2_P4_datai )) ;8253
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8254");		//(= P2_P4_addr    P2_P4_tail )) ;8254
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8255");		//(= P2_P4_rd    0b1)) ;8255
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8256");		//(= P2_P4_mf    0b10)) ;8256
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8257");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8257
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8258");		//(= P2_P4_rd    0b1)) ;8258
                                                                P2_P4_m = P2_P4_datai; $display(";A 8259");		//(= P2_P4_m    P2_P4_datai )) ;8259
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8260");		//(= P2_P4_mf    0b11)) ;8260
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8261");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8261
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8262");		//(= P2_P4_rd    0b1)) ;8262
                                                                P2_P4_m = P2_P4_datai; $display(";A 8263");		//(= P2_P4_m    P2_P4_datai )) ;8263
                                                            end
                                                    endcase
                                                    P2_P4_t = 32'sb00000000000000000000000000000000; $display(";A 8264");		//(= P2_P4_t    0b00000000000000000000000000000000)) ;8264
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8265");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8265
                                                                P2_P4_reg0 = (P2_P4_t - P2_P4_m); $display(";A 8266");		//(= P2_P4_reg0    (bv-sub P2_P4_t  P2_P4_m ))) ;8266
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8267");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8267
                                                                P2_P4_reg1 = (P2_P4_t - P2_P4_m); $display(";A 8268");		//(= P2_P4_reg1    (bv-sub P2_P4_t  P2_P4_m ))) ;8268
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8269");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8269
                                                                P2_P4_reg2 = (P2_P4_t - P2_P4_m); $display(";A 8270");		//(= P2_P4_reg2    (bv-sub P2_P4_t  P2_P4_m ))) ;8270
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8271");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8271
                                                                P2_P4_reg3 = (P2_P4_t - P2_P4_m); $display(";A 8272");		//(= P2_P4_reg3    (bv-sub P2_P4_t  P2_P4_m ))) ;8272
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8273");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8273
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0001 :
                                                begin
                                                    $display(";A 8274");		//(= P2_P4_ff    0b0001)) ;8274
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8275");		//(= P2_P4_mf    0b00)) ;8275
                                                                P2_P4_m = P2_P4_tail; $display(";A 8276");		//(= P2_P4_m    P2_P4_tail )) ;8276
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8277");		//(= P2_P4_mf    0b01)) ;8277
                                                                P2_P4_m = P2_P4_datai; $display(";A 8278");		//(= P2_P4_m    P2_P4_datai )) ;8278
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8279");		//(= P2_P4_addr    P2_P4_tail )) ;8279
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8280");		//(= P2_P4_rd    0b1)) ;8280
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8281");		//(= P2_P4_mf    0b10)) ;8281
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8282");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8282
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8283");		//(= P2_P4_rd    0b1)) ;8283
                                                                P2_P4_m = P2_P4_datai; $display(";A 8284");		//(= P2_P4_m    P2_P4_datai )) ;8284
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8285");		//(= P2_P4_mf    0b11)) ;8285
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8286");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8286
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8287");		//(= P2_P4_rd    0b1)) ;8287
                                                                P2_P4_m = P2_P4_datai; $display(";A 8288");		//(= P2_P4_m    P2_P4_datai )) ;8288
                                                            end
                                                    endcase
                                                    P2_P4_reg2 = P2_P4_reg3; $display(";A 8289");		//(= P2_P4_reg2    P2_P4_reg3 )) ;8289
                                                    P2_P4_reg3 = P2_P4_m; $display(";A 8290");		//(= P2_P4_reg3    P2_P4_m )) ;8290
                                                end
                                            4'b0010 :
                                                begin
                                                    $display(";A 8291");		//(= P2_P4_ff    0b0010)) ;8291
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8292");		//(= P2_P4_mf    0b00)) ;8292
                                                                P2_P4_m = P2_P4_tail; $display(";A 8293");		//(= P2_P4_m    P2_P4_tail )) ;8293
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8294");		//(= P2_P4_mf    0b01)) ;8294
                                                                P2_P4_m = P2_P4_datai; $display(";A 8295");		//(= P2_P4_m    P2_P4_datai )) ;8295
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8296");		//(= P2_P4_addr    P2_P4_tail )) ;8296
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8297");		//(= P2_P4_rd    0b1)) ;8297
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8298");		//(= P2_P4_mf    0b10)) ;8298
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8299");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8299
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8300");		//(= P2_P4_rd    0b1)) ;8300
                                                                P2_P4_m = P2_P4_datai; $display(";A 8301");		//(= P2_P4_m    P2_P4_datai )) ;8301
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8302");		//(= P2_P4_mf    0b11)) ;8302
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8303");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8303
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8304");		//(= P2_P4_rd    0b1)) ;8304
                                                                P2_P4_m = P2_P4_datai; $display(";A 8305");		//(= P2_P4_m    P2_P4_datai )) ;8305
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8306");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8306
                                                                P2_P4_reg0 = P2_P4_m; $display(";A 8307");		//(= P2_P4_reg0    P2_P4_m )) ;8307
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8308");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8308
                                                                P2_P4_reg1 = P2_P4_m; $display(";A 8309");		//(= P2_P4_reg1    P2_P4_m )) ;8309
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8310");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8310
                                                                P2_P4_reg2 = P2_P4_m; $display(";A 8311");		//(= P2_P4_reg2    P2_P4_m )) ;8311
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8312");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8312
                                                                P2_P4_reg3 = P2_P4_m; $display(";A 8313");		//(= P2_P4_reg3    P2_P4_m )) ;8313
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8314");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8314
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0011 :
                                                begin
                                                    $display(";A 8315");		//(= P2_P4_ff    0b0011)) ;8315
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8316");		//(= P2_P4_mf    0b00)) ;8316
                                                                P2_P4_m = P2_P4_tail; $display(";A 8317");		//(= P2_P4_m    P2_P4_tail )) ;8317
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8318");		//(= P2_P4_mf    0b01)) ;8318
                                                                P2_P4_m = P2_P4_datai; $display(";A 8319");		//(= P2_P4_m    P2_P4_datai )) ;8319
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8320");		//(= P2_P4_addr    P2_P4_tail )) ;8320
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8321");		//(= P2_P4_rd    0b1)) ;8321
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8322");		//(= P2_P4_mf    0b10)) ;8322
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8323");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8323
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8324");		//(= P2_P4_rd    0b1)) ;8324
                                                                P2_P4_m = P2_P4_datai; $display(";A 8325");		//(= P2_P4_m    P2_P4_datai )) ;8325
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8326");		//(= P2_P4_mf    0b11)) ;8326
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8327");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8327
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8328");		//(= P2_P4_rd    0b1)) ;8328
                                                                P2_P4_m = P2_P4_datai; $display(";A 8329");		//(= P2_P4_m    P2_P4_datai )) ;8329
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8330");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8330
                                                                P2_P4_reg0 = P2_P4_m; $display(";A 8331");		//(= P2_P4_reg0    P2_P4_m )) ;8331
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8332");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8332
                                                                P2_P4_reg1 = P2_P4_m; $display(";A 8333");		//(= P2_P4_reg1    P2_P4_m )) ;8333
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8334");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8334
                                                                P2_P4_reg2 = P2_P4_m; $display(";A 8335");		//(= P2_P4_reg2    P2_P4_m )) ;8335
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8336");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8336
                                                                P2_P4_reg3 = P2_P4_m; $display(";A 8337");		//(= P2_P4_reg3    P2_P4_m )) ;8337
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8338");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8338
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0100 :
                                                begin
                                                    $display(";A 8339");		//(= P2_P4_ff    0b0100)) ;8339
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8340");		//(= P2_P4_mf    0b00)) ;8340
                                                                P2_P4_m = P2_P4_tail; $display(";A 8341");		//(= P2_P4_m    P2_P4_tail )) ;8341
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8342");		//(= P2_P4_mf    0b01)) ;8342
                                                                P2_P4_m = P2_P4_datai; $display(";A 8343");		//(= P2_P4_m    P2_P4_datai )) ;8343
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8344");		//(= P2_P4_addr    P2_P4_tail )) ;8344
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8345");		//(= P2_P4_rd    0b1)) ;8345
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8346");		//(= P2_P4_mf    0b10)) ;8346
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8347");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8347
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8348");		//(= P2_P4_rd    0b1)) ;8348
                                                                P2_P4_m = P2_P4_datai; $display(";A 8349");		//(= P2_P4_m    P2_P4_datai )) ;8349
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8350");		//(= P2_P4_mf    0b11)) ;8350
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8351");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8351
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8352");		//(= P2_P4_rd    0b1)) ;8352
                                                                P2_P4_m = P2_P4_datai; $display(";A 8353");		//(= P2_P4_m    P2_P4_datai )) ;8353
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8354");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8354
                                                                P2_P4_reg0 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8355");		//(= P2_P4_reg0    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8355
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8356");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8356
                                                                P2_P4_reg1 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8357");		//(= P2_P4_reg1    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8357
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8358");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8358
                                                                P2_P4_reg2 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8359");		//(= P2_P4_reg2    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8359
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8360");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8360
                                                                P2_P4_reg3 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8361");		//(= P2_P4_reg3    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8361
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8362");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8362
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0101 :
                                                begin
                                                    $display(";A 8363");		//(= P2_P4_ff    0b0101)) ;8363
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8364");		//(= P2_P4_mf    0b00)) ;8364
                                                                P2_P4_m = P2_P4_tail; $display(";A 8365");		//(= P2_P4_m    P2_P4_tail )) ;8365
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8366");		//(= P2_P4_mf    0b01)) ;8366
                                                                P2_P4_m = P2_P4_datai; $display(";A 8367");		//(= P2_P4_m    P2_P4_datai )) ;8367
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8368");		//(= P2_P4_addr    P2_P4_tail )) ;8368
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8369");		//(= P2_P4_rd    0b1)) ;8369
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8370");		//(= P2_P4_mf    0b10)) ;8370
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8371");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8371
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8372");		//(= P2_P4_rd    0b1)) ;8372
                                                                P2_P4_m = P2_P4_datai; $display(";A 8373");		//(= P2_P4_m    P2_P4_datai )) ;8373
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8374");		//(= P2_P4_mf    0b11)) ;8374
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8375");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8375
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8376");		//(= P2_P4_rd    0b1)) ;8376
                                                                P2_P4_m = P2_P4_datai; $display(";A 8377");		//(= P2_P4_m    P2_P4_datai )) ;8377
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8378");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8378
                                                                P2_P4_reg0 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8379");		//(= P2_P4_reg0    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8379
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8380");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8380
                                                                P2_P4_reg1 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8381");		//(= P2_P4_reg1    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8381
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8382");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8382
                                                                P2_P4_reg2 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8383");		//(= P2_P4_reg2    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8383
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8384");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8384
                                                                P2_P4_reg3 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8385");		//(= P2_P4_reg3    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8385
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8386");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8386
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0110 :
                                                begin
                                                    $display(";A 8387");		//(= P2_P4_ff    0b0110)) ;8387
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8388");		//(= P2_P4_mf    0b00)) ;8388
                                                                P2_P4_m = P2_P4_tail; $display(";A 8389");		//(= P2_P4_m    P2_P4_tail )) ;8389
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8390");		//(= P2_P4_mf    0b01)) ;8390
                                                                P2_P4_m = P2_P4_datai; $display(";A 8391");		//(= P2_P4_m    P2_P4_datai )) ;8391
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8392");		//(= P2_P4_addr    P2_P4_tail )) ;8392
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8393");		//(= P2_P4_rd    0b1)) ;8393
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8394");		//(= P2_P4_mf    0b10)) ;8394
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8395");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8395
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8396");		//(= P2_P4_rd    0b1)) ;8396
                                                                P2_P4_m = P2_P4_datai; $display(";A 8397");		//(= P2_P4_m    P2_P4_datai )) ;8397
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8398");		//(= P2_P4_mf    0b11)) ;8398
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8399");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8399
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8400");		//(= P2_P4_rd    0b1)) ;8400
                                                                P2_P4_m = P2_P4_datai; $display(";A 8401");		//(= P2_P4_m    P2_P4_datai )) ;8401
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8402");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8402
                                                                P2_P4_reg0 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8403");		//(= P2_P4_reg0    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8403
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8404");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8404
                                                                P2_P4_reg1 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8405");		//(= P2_P4_reg1    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8405
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8406");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8406
                                                                P2_P4_reg2 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8407");		//(= P2_P4_reg2    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8407
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8408");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8408
                                                                P2_P4_reg3 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8409");		//(= P2_P4_reg3    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8409
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8410");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8410
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b0111 :
                                                begin
                                                    $display(";A 8411");		//(= P2_P4_ff    0b0111)) ;8411
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8412");		//(= P2_P4_mf    0b00)) ;8412
                                                                P2_P4_m = P2_P4_tail; $display(";A 8413");		//(= P2_P4_m    P2_P4_tail )) ;8413
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8414");		//(= P2_P4_mf    0b01)) ;8414
                                                                P2_P4_m = P2_P4_datai; $display(";A 8415");		//(= P2_P4_m    P2_P4_datai )) ;8415
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8416");		//(= P2_P4_addr    P2_P4_tail )) ;8416
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8417");		//(= P2_P4_rd    0b1)) ;8417
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8418");		//(= P2_P4_mf    0b10)) ;8418
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8419");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8419
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8420");		//(= P2_P4_rd    0b1)) ;8420
                                                                P2_P4_m = P2_P4_datai; $display(";A 8421");		//(= P2_P4_m    P2_P4_datai )) ;8421
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8422");		//(= P2_P4_mf    0b11)) ;8422
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8423");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8423
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8424");		//(= P2_P4_rd    0b1)) ;8424
                                                                P2_P4_m = P2_P4_datai; $display(";A 8425");		//(= P2_P4_m    P2_P4_datai )) ;8425
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8426");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8426
                                                                P2_P4_reg0 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8427");		//(= P2_P4_reg0    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8427
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8428");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8428
                                                                P2_P4_reg1 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8429");		//(= P2_P4_reg1    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8429
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8430");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8430
                                                                P2_P4_reg2 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8431");		//(= P2_P4_reg2    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8431
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8432");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8432
                                                                P2_P4_reg3 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8433");		//(= P2_P4_reg3    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8433
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8434");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8434
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1000 :
                                                begin
                                                    $display(";A 8435");		//(= P2_P4_ff    0b1000)) ;8435
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8436");		//(= P2_P4_mf    0b00)) ;8436
                                                                P2_P4_m = P2_P4_tail; $display(";A 8437");		//(= P2_P4_m    P2_P4_tail )) ;8437
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8438");		//(= P2_P4_mf    0b01)) ;8438
                                                                P2_P4_m = P2_P4_datai; $display(";A 8439");		//(= P2_P4_m    P2_P4_datai )) ;8439
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8440");		//(= P2_P4_addr    P2_P4_tail )) ;8440
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8441");		//(= P2_P4_rd    0b1)) ;8441
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8442");		//(= P2_P4_mf    0b10)) ;8442
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8443");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8443
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8444");		//(= P2_P4_rd    0b1)) ;8444
                                                                P2_P4_m = P2_P4_datai; $display(";A 8445");		//(= P2_P4_m    P2_P4_datai )) ;8445
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8446");		//(= P2_P4_mf    0b11)) ;8446
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8447");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8447
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8448");		//(= P2_P4_rd    0b1)) ;8448
                                                                P2_P4_m = P2_P4_datai; $display(";A 8449");		//(= P2_P4_m    P2_P4_datai )) ;8449
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8450");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8450
                                                                P2_P4_reg0 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8451");		//(= P2_P4_reg0    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8451
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8452");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8452
                                                                P2_P4_reg1 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8453");		//(= P2_P4_reg1    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8453
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8454");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8454
                                                                P2_P4_reg2 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8455");		//(= P2_P4_reg2    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8455
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8456");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8456
                                                                P2_P4_reg3 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8457");		//(= P2_P4_reg3    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8457
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8458");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8458
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1001 :
                                                begin
                                                    $display(";A 8459");		//(= P2_P4_ff    0b1001)) ;8459
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8460");		//(= P2_P4_mf    0b00)) ;8460
                                                                P2_P4_m = P2_P4_tail; $display(";A 8461");		//(= P2_P4_m    P2_P4_tail )) ;8461
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8462");		//(= P2_P4_mf    0b01)) ;8462
                                                                P2_P4_m = P2_P4_datai; $display(";A 8463");		//(= P2_P4_m    P2_P4_datai )) ;8463
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8464");		//(= P2_P4_addr    P2_P4_tail )) ;8464
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8465");		//(= P2_P4_rd    0b1)) ;8465
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8466");		//(= P2_P4_mf    0b10)) ;8466
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8467");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8467
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8468");		//(= P2_P4_rd    0b1)) ;8468
                                                                P2_P4_m = P2_P4_datai; $display(";A 8469");		//(= P2_P4_m    P2_P4_datai )) ;8469
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8470");		//(= P2_P4_mf    0b11)) ;8470
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8471");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8471
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8472");		//(= P2_P4_rd    0b1)) ;8472
                                                                P2_P4_m = P2_P4_datai; $display(";A 8473");		//(= P2_P4_m    P2_P4_datai )) ;8473
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8474");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8474
                                                                P2_P4_reg0 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8475");		//(= P2_P4_reg0    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8475
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8476");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8476
                                                                P2_P4_reg1 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8477");		//(= P2_P4_reg1    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8477
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8478");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8478
                                                                P2_P4_reg2 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8479");		//(= P2_P4_reg2    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8479
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8480");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8480
                                                                P2_P4_reg3 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8481");		//(= P2_P4_reg3    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8481
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8482");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8482
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1010 :
                                                begin
                                                    $display(";A 8483");		//(= P2_P4_ff    0b1010)) ;8483
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8484");		//(= P2_P4_mf    0b00)) ;8484
                                                                P2_P4_m = P2_P4_tail; $display(";A 8485");		//(= P2_P4_m    P2_P4_tail )) ;8485
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8486");		//(= P2_P4_mf    0b01)) ;8486
                                                                P2_P4_m = P2_P4_datai; $display(";A 8487");		//(= P2_P4_m    P2_P4_datai )) ;8487
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8488");		//(= P2_P4_addr    P2_P4_tail )) ;8488
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8489");		//(= P2_P4_rd    0b1)) ;8489
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8490");		//(= P2_P4_mf    0b10)) ;8490
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8491");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8491
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8492");		//(= P2_P4_rd    0b1)) ;8492
                                                                P2_P4_m = P2_P4_datai; $display(";A 8493");		//(= P2_P4_m    P2_P4_datai )) ;8493
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8494");		//(= P2_P4_mf    0b11)) ;8494
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8495");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8495
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8496");		//(= P2_P4_rd    0b1)) ;8496
                                                                P2_P4_m = P2_P4_datai; $display(";A 8497");		//(= P2_P4_m    P2_P4_datai )) ;8497
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8498");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8498
                                                                P2_P4_reg0 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8499");		//(= P2_P4_reg0    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8499
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8500");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8500
                                                                P2_P4_reg1 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8501");		//(= P2_P4_reg1    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8501
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8502");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8502
                                                                P2_P4_reg2 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8503");		//(= P2_P4_reg2    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8503
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8504");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8504
                                                                P2_P4_reg3 = ((P2_P4_r + P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8505");		//(= P2_P4_reg3    (bv-smod (bv-add P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8505
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8506");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8506
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1011 :
                                                begin
                                                    $display(";A 8507");		//(= P2_P4_ff    0b1011)) ;8507
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8508");		//(= P2_P4_mf    0b00)) ;8508
                                                                P2_P4_m = P2_P4_tail; $display(";A 8509");		//(= P2_P4_m    P2_P4_tail )) ;8509
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8510");		//(= P2_P4_mf    0b01)) ;8510
                                                                P2_P4_m = P2_P4_datai; $display(";A 8511");		//(= P2_P4_m    P2_P4_datai )) ;8511
                                                                P2_P4_addr <= #1 P2_P4_tail; $display(";A 8512");		//(= P2_P4_addr    P2_P4_tail )) ;8512
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8513");		//(= P2_P4_rd    0b1)) ;8513
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8514");		//(= P2_P4_mf    0b10)) ;8514
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg1) % 32'b00000000000100000000000000000000); $display(";A 8515");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg1 ) 0b00000000000100000000000000000000))) ;8515
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8516");		//(= P2_P4_rd    0b1)) ;8516
                                                                P2_P4_m = P2_P4_datai; $display(";A 8517");		//(= P2_P4_m    P2_P4_datai )) ;8517
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8518");		//(= P2_P4_mf    0b11)) ;8518
                                                                P2_P4_addr <= #1 ((P2_P4_tail + P2_P4_reg2) % 32'b00000000000100000000000000000000); $display(";A 8519");		//(= P2_P4_addr    (bv-smod (bv-add P2_P4_tail  P2_P4_reg2 ) 0b00000000000100000000000000000000))) ;8519
                                                                P2_P4_rd <= #1 1'b1; $display(";A 8520");		//(= P2_P4_rd    0b1)) ;8520
                                                                P2_P4_m = P2_P4_datai; $display(";A 8521");		//(= P2_P4_m    P2_P4_datai )) ;8521
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8522");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8522
                                                                P2_P4_reg0 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8523");		//(= P2_P4_reg0    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8523
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8524");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8524
                                                                P2_P4_reg1 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8525");		//(= P2_P4_reg1    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8525
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8526");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8526
                                                                P2_P4_reg2 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8527");		//(= P2_P4_reg2    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8527
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8528");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8528
                                                                P2_P4_reg3 = ((P2_P4_r - P2_P4_m) % 32'b00000000000000000000000000000000); $display(";A 8529");		//(= P2_P4_reg3    (bv-smod (bv-sub P2_P4_r  P2_P4_m ) 0b00000000000000000000000000000000))) ;8529
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8530");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8530
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1100 :
                                                begin
                                                    $display(";A 8531");		//(= P2_P4_ff    0b1100)) ;8531
                                                    case (P2_P4_mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 8532");		//(= P2_P4_mf    0b00)) ;8532
                                                                P2_P4_t = (P2_P4_r / 32'sb00000000000000000000000000000010); $display(";A 8533");		//(= P2_P4_t    (bv-sdiv P2_P4_r  0b00000000000000000000000000000010))) ;8533
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 8534");		//(= P2_P4_mf    0b01)) ;8534
                                                                P2_P4_t = (P2_P4_r / 32'sb00000000000000000000000000000010); $display(";A 8535");		//(= P2_P4_t    (bv-sdiv P2_P4_r  0b00000000000000000000000000000010))) ;8535
                                                                if ((P2_P4_B == 1'b1)) begin
                                                                    $display(";A 8536");		//(= (bv-comp P2_P4_B  0b1)   0b1)) ;8536
                                                                    P2_P4_t = (P2_P4_t % 32'b00100000000000000000000000000000); $display(";A 8538");		//(= P2_P4_t    (bv-smod P2_P4_t  0b00100000000000000000000000000000))) ;8538
                                                                end
                                                                else begin
                                                                    $display(";A 8537");		//(= (bv-comp P2_P4_B  0b1)   0b0)) ;8537
                                                                end
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 8539");		//(= P2_P4_mf    0b10)) ;8539
                                                                P2_P4_t = ((P2_P4_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 8540");		//(= P2_P4_t    (bv-mul (bv-smod P2_P4_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;8540
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 8541");		//(= P2_P4_mf    0b11)) ;8541
                                                                P2_P4_t = ((P2_P4_r % 32'b00100000000000000000000000000000) * 32'b00000000000000000000000000000010); $display(";A 8542");		//(= P2_P4_t    (bv-mul (bv-smod P2_P4_r  0b00100000000000000000000000000000) 0b00000000000000000000000000000010))) ;8542
                                                                if ((P2_P4_t > 32'b11111111111111111111111111111111)) begin
                                                                    $display(";A 8543");		//(= (bool-to-bv (bv-gt P2_P4_t  0b11111111111111111111111111111111))   0b1)) ;8543
                                                                    P2_P4_B = 1'b1; $display(";A 8545");		//(= P2_P4_B    0b1)) ;8545
                                                                end
                                                                else begin
                                                                    $display(";A 8544");		//(= (bool-to-bv (bv-gt P2_P4_t  0b11111111111111111111111111111111))   0b0)) ;8544
                                                                    P2_P4_B = 1'b0; $display(";A 8546");		//(= P2_P4_B    0b0)) ;8546
                                                                end
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8547");		//(= (and (/= P2_P4_mf  0b00) (/= P2_P4_mf  0b01) (/= P2_P4_mf  0b10) (/= P2_P4_mf  0b11))   true)) ;8547
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                    case (P2_P4_d)
                                                        32'sb00000000000000000000000000000000 :
                                                            begin
                                                                $display(";A 8548");		//(= P2_P4_d    0b00000000000000000000000000000000)) ;8548
                                                                P2_P4_reg0 = P2_P4_t; $display(";A 8549");		//(= P2_P4_reg0    P2_P4_t )) ;8549
                                                            end
                                                        32'sb00000000000000000000000000000001 :
                                                            begin
                                                                $display(";A 8550");		//(= P2_P4_d    0b00000000000000000000000000000001)) ;8550
                                                                P2_P4_reg1 = P2_P4_t; $display(";A 8551");		//(= P2_P4_reg1    P2_P4_t )) ;8551
                                                            end
                                                        32'sb00000000000000000000000000000010 :
                                                            begin
                                                                $display(";A 8552");		//(= P2_P4_d    0b00000000000000000000000000000010)) ;8552
                                                                P2_P4_reg2 = P2_P4_t; $display(";A 8553");		//(= P2_P4_reg2    P2_P4_t )) ;8553
                                                            end
                                                        32'sb00000000000000000000000000000011 :
                                                            begin
                                                                $display(";A 8554");		//(= P2_P4_d    0b00000000000000000000000000000011)) ;8554
                                                                P2_P4_reg3 = P2_P4_t; $display(";A 8555");		//(= P2_P4_reg3    P2_P4_t )) ;8555
                                                            end
                                                        default:
                                                            begin
                                                                $display(";A 8556");		//(= (and (/= P2_P4_d  0b00000000000000000000000000000000) (/= P2_P4_d  0b00000000000000000000000000000001) (/= P2_P4_d  0b00000000000000000000000000000010) (/= P2_P4_d  0b00000000000000000000000000000011))   true)) ;8556
                                                                begin
                                                                end
                                                            end
                                                    endcase
                                                end
                                            4'b1101 :
                                                begin
                                                    $display(";A 8557");		//(= P2_P4_ff    0b1101)) ;8557
                                                    begin
                                                    end
                                                end
                                            4'b1110 :
                                                begin
                                                    $display(";A 8558");		//(= P2_P4_ff    0b1110)) ;8558
                                                    begin
                                                    end
                                                end
                                            4'b1111 :
                                                begin
                                                    $display(";A 8559");		//(= P2_P4_ff    0b1111)) ;8559
                                                    begin
                                                    end
                                                end
                                        endcase
                                    end
                                    else begin
                                        $display(";A 8226");		//(= (bv-not (bv-comp P2_P4_df  0b00000000000000000000000000000111))   0b0)) ;8226
                                        if ((P2_P4_df == 32'b00000000000000000000000000000111)) begin
                                            $display(";A 8560");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000111)   0b1)) ;8560
                                            case (P2_P4_mf)
                                                2'b00 :
                                                    begin
                                                        $display(";A 8562");		//(= P2_P4_mf    0b00)) ;8562
                                                        P2_P4_m = P2_P4_tail; $display(";A 8563");		//(= P2_P4_m    P2_P4_tail )) ;8563
                                                    end
                                                2'b01 :
                                                    begin
                                                        $display(";A 8564");		//(= P2_P4_mf    0b01)) ;8564
                                                        P2_P4_m = P2_P4_tail; $display(";A 8565");		//(= P2_P4_m    P2_P4_tail )) ;8565
                                                    end
                                                2'b10 :
                                                    begin
                                                        $display(";A 8566");		//(= P2_P4_mf    0b10)) ;8566
                                                        P2_P4_m = ((P2_P4_reg1 % 32'b00000000000100000000000000000000) + (P2_P4_tail % 32'b00000000000100000000000000000000)); $display(";A 8567");		//(= P2_P4_m    (bv-add (bv-smod P2_P4_reg1  0b00000000000100000000000000000000) (bv-smod P2_P4_tail  0b00000000000100000000000000000000)))) ;8567
                                                    end
                                                2'b11 :
                                                    begin
                                                        $display(";A 8568");		//(= P2_P4_mf    0b11)) ;8568
                                                        P2_P4_m = ((P2_P4_reg2 % 32'b00000000000100000000000000000000) + (P2_P4_tail % 32'b00000000000100000000000000000000)); $display(";A 8569");		//(= P2_P4_m    (bv-add (bv-smod P2_P4_reg2  0b00000000000100000000000000000000) (bv-smod P2_P4_tail  0b00000000000100000000000000000000)))) ;8569
                                                    end
                                            endcase
                                            P2_P4_addr <= #1 ((P2_P4_m % 32'sb00000000000000000000000000000010) * 32'sb00000000000000000000000000010100); $display(";A 8570");		//(= P2_P4_addr    (bv-mul (bv-smod P2_P4_m  0b00000000000000000000000000000010) 0b00000000000000000000000000010100))) ;8570
                                            P2_P4_wr <= #1 1'b1; $display(";A 8571");		//(= P2_P4_wr    0b1)) ;8571
                                            P2_P4_datao <= #1 P2_P4_r; $display(";A 8572");		//(= P2_P4_datao    P2_P4_r )) ;8572
                                        end
                                        else begin
                                            $display(";A 8561");		//(= (bv-comp P2_P4_df  0b00000000000000000000000000000111)   0b0)) ;8561
                                        end
                                    end
                                end
                        endcase
                        P2_P4_state = 1'sb0; $display(";A 8573");		//(= P2_P4_state    0b0)) ;8573
                    end
            endcase
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:13072
    always @(P2_td2 or P2_td1 or P2_din or P2_sel or P2_tad4 or P2_tad3 or P2_ad22 or P2_ad21 or P2_ad12 or P2_ad11 or P2_do4 or P2_do3 or P2_tad1 or P2_ad41 or P2_wr4 or P2_tad2 or P2_ad31 or P2_wr3 or P2_as11 or P2_as21 or P2_as22 or P2_dc2 or P2_mio2 or P2_wr2 or P2_rd4 or P2_do2 or P2_as12 or P2_dc1 or P2_mio1 or P2_wr1 or P2_rd3 or P2_do1) begin
        P2_di3 <= #1 (P2_do1 % 32'b00000000000100000000000000000000); $display(";A 8574");		//(= P2_di3    (bv-smod P2_do1  0b00000000000100000000000000000000))) ;8574
        P2_r12 <= #1 (~((((P2_rd3 & P2_wr1) & P2_mio1) & P2_dc1) & (~P2_as12))); $display(";A 8575");		//(= P2_r12    (bv-not (bv-and (bv-and (bv-and (bv-and P2_rd3  P2_wr1 ) P2_mio1 ) P2_dc1 ) (bv-not P2_as12 ))))) ;8575
        P2_di4 <= #1 P2_do2; $display(";A 8576");		//(= P2_di4    P2_do2 )) ;8576
        P2_r22 <= #1 (~((((P2_rd4 & P2_wr2) & P2_mio2) & P2_dc2) & (~P2_as22))); $display(";A 8577");		//(= P2_r22    (bv-not (bv-and (bv-and (bv-and (bv-and P2_rd4  P2_wr2 ) P2_mio2 ) P2_dc2 ) (bv-not P2_as22 ))))) ;8577
        P2_r11 <= #1 P2_as21; $display(";A 8578");		//(= P2_r11    P2_as21 )) ;8578
        P2_r21 <= #1 P2_as11; $display(";A 8579");		//(= P2_r21    P2_as11 )) ;8579
        if ((P2_wr3 == 1'b1)) begin
            $display(";A 8580");		//(= (bv-comp P2_wr3  0b1)   0b1)) ;8580
            P2_tad3 <= #1 P2_ad31; $display(";A 8582");		//(= P2_tad3    P2_ad31 )) ;8582
        end
        else begin
            $display(";A 8581");		//(= (bv-comp P2_wr3  0b1)   0b0)) ;8581
            P2_tad3 <= #1 (P2_tad2 % 30'b000000000100000000000000000000); $display(";A 8583");		//(= P2_tad3    (bv-smod P2_tad2  0b000000000100000000000000000000))) ;8583
        end
        if ((P2_wr4 == 1'b1)) begin
            $display(";A 8584");		//(= (bv-comp P2_wr4  0b1)   0b1)) ;8584
            P2_tad4 <= #1 P2_ad41; $display(";A 8586");		//(= P2_tad4    P2_ad41 )) ;8586
        end
        else begin
            $display(";A 8585");		//(= (bv-comp P2_wr4  0b1)   0b0)) ;8585
            P2_tad4 <= #1 (P2_tad1 % 30'b000000000100000000000000000000); $display(";A 8587");		//(= P2_tad4    (bv-smod P2_tad1  0b000000000100000000000000000000))) ;8587
        end
        if ((P2_do3 > 32'b00010000000000000000000000000000)) begin
            $display(";A 8588");		//(= (bool-to-bv (bv-gt P2_do3  0b00010000000000000000000000000000))   0b1)) ;8588
            P2_tad1 <= #1 P2_ad11; $display(";A 8590");		//(= P2_tad1    P2_ad11 )) ;8590
        end
        else begin
            $display(";A 8589");		//(= (bool-to-bv (bv-gt P2_do3  0b00010000000000000000000000000000))   0b0)) ;8589
            P2_tad1 <= #1 P2_ad12; $display(";A 8591");		//(= P2_tad1    P2_ad12 )) ;8591
        end
        if ((P2_do4 > 32'b00100000000000000000000000000000)) begin
            $display(";A 8592");		//(= (bool-to-bv (bv-gt P2_do4  0b00100000000000000000000000000000))   0b1)) ;8592
            P2_tad2 <= #1 P2_ad21; $display(";A 8594");		//(= P2_tad2    P2_ad21 )) ;8594
        end
        else begin
            $display(";A 8593");		//(= (bool-to-bv (bv-gt P2_do4  0b00100000000000000000000000000000))   0b0)) ;8593
            P2_tad2 <= #1 P2_ad22; $display(";A 8595");		//(= P2_tad2    P2_ad22 )) ;8595
        end
        P2_dout <= #1 ((P2_tad3 * P2_tad4) % 20'b10000000000000000000); $display(";A 8596");		//(= P2_dout    (bv-smod (bv-mul P2_tad3  P2_tad4 ) 0b10000000000000000000))) ;8596
        if ((P2_sel == 1'b0)) begin
            $display(";A 8597");		//(= (bv-comp P2_sel  0b0)   0b1)) ;8597
            P2_td1 <= #1 32'sb00000000000000000000000000000000; $display(";A 8599");		//(= P2_td1    0b00000000000000000000000000000000)) ;8599
            P2_td2 <= #1 P2_din; $display(";A 8600");		//(= P2_td2    P2_din )) ;8600
        end
        else begin
            $display(";A 8598");		//(= (bv-comp P2_sel  0b0)   0b0)) ;8598
            P2_td1 <= #1 P2_din; $display(";A 8601");		//(= P2_td1    P2_din )) ;8601
            P2_td2 <= #1 32'sb00000000000000000000000000000000; $display(";A 8602");		//(= P2_td2    0b00000000000000000000000000000000)) ;8602
        end
        P2_di1 <= #1 (P2_do4 * P2_td1); $display(";A 8603");		//(= P2_di1    (bv-mul P2_do4  P2_td1 ))) ;8603
        P2_di2 <= #1 (P2_do3 * P2_td2); $display(";A 8604");		//(= P2_di2    (bv-mul P2_do3  P2_td2 ))) ;8604
        P2_aux <= #1 ((P2_tad1 * P2_tad2) % 30'b000000000000000000000000001000); $display(";A 8605");		//(= P2_aux    (bv-smod (bv-mul P2_tad1  P2_tad2 ) 0b000000000000000000000000001000))) ;8605
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:13113
    always @(posedge reset or posedge clock) begin
        if ((reset == 1'b1)) begin
            sel1 <= #1 1'b0; $display(";A 8608");		//(= sel1    0b0)) ;8608
            sel2 <= #1 1'b0; $display(";A 8609");		//(= sel2    0b0)) ;8609
        end
        else begin
            if ((do1 == 32'b00000000000000000000000000100111)) begin
                $display(";A 8610");		//(= (bv-comp do1  0b00000000000000000000000000100111)   0b1)) ;8610
                sel2 <= #1 1'b1; $display(";A 8612");		//(= sel2    0b1)) ;8612
            end
            else begin
                $display(";A 8611");		//(= (bv-comp do1  0b00000000000000000000000000100111)   0b0)) ;8611
                if ((do1 == 32'b00000000000000000000011011000111)) begin
                    $display(";A 8613");		//(= (bv-comp do1  0b00000000000000000000011011000111)   0b1)) ;8613
                    sel2 <= #1 1'b0; $display(";A 8615");		//(= sel2    0b0)) ;8615
                end
                else begin
                    $display(";A 8614");		//(= (bv-comp do1  0b00000000000000000000011011000111)   0b0)) ;8614
                end
            end
            if ((do2 == 32'b00000000000000000000000110001110)) begin
                $display(";A 8616");		//(= (bv-comp do2  0b00000000000000000000000110001110)   0b1)) ;8616
                sel1 <= #1 1'b1; $display(";A 8618");		//(= sel1    0b1)) ;8618
            end
            else begin
                $display(";A 8617");		//(= (bv-comp do2  0b00000000000000000000000110001110)   0b0)) ;8617
                if ((do2 == 32'b00000000000000000000001111110101)) begin
                    $display(";A 8619");		//(= (bv-comp do2  0b00000000000000000000001111110101)   0b1)) ;8619
                    sel1 <= #1 1'b0; $display(";A 8621");		//(= sel1    0b0)) ;8621
                end
                else begin
                    $display(";A 8620");		//(= (bv-comp do2  0b00000000000000000000001111110101)   0b0)) ;8620
                end
            end
        end
    end

    // Following code segment is generated from /home/ziyue/researchlib/Micro_Eletronic/STSearch/tests/b19/src/b19.v:13133
    always @(ax2 or ax1 or do2 or do1 or in3 or in2 or in1 or sel2 or sel1) begin
        if (((sel1 == 1'b0) & (sel2 == 1'b1))) begin
            $display(";A 8622");		//(= (bv-and (bv-comp sel1  0b0) (bv-comp sel2  0b1))   0b1)) ;8622
            di1 <= #1 (in1 / 32'b00000000000000000000000000000010); $display(";A 8624");		//(= di1    (bv-sdiv in1  0b00000000000000000000000000000010))) ;8624
            di2 <= #1 (in2 / 32'b00000000000000000000000000010000); $display(";A 8625");		//(= di2    (bv-sdiv in2  0b00000000000000000000000000010000))) ;8625
        end
        else begin
            $display(";A 8623");		//(= (bv-and (bv-comp sel1  0b0) (bv-comp sel2  0b1))   0b0)) ;8623
            di1 <= #1 (in1 / 32'b00000000000000000000000000000010); $display(";A 8626");		//(= di1    (bv-sdiv in1  0b00000000000000000000000000000010))) ;8626
            di2 <= #1 (in2 / 32'b00000000000000000000000000001000); $display(";A 8627");		//(= di2    (bv-sdiv in2  0b00000000000000000000000000001000))) ;8627
        end
        ris <= #1 (((ax1 - ax2) * do1) - ((ax1 - ax2) * do2)); $display(";A 8628");		//(= ris    (bv-sub (bv-mul (bv-sub ax1  ax2 ) do1 ) (bv-mul (bv-sub ax1  ax2 ) do2 )))) ;8628
    end

endmodule

