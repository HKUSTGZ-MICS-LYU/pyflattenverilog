
	//`define CODE_FOR_SYNTHESIS				// uncomment this macro will remove all non-systhesis code
	`define USE_SIMULATION_CODE					// uncomment this to use simulation instruction memory
	
	`define PC_WIDTH				8
	`define	INSTR_MEM_ADDR_WIDTH	8
	`define DATA_MEM_ADDR_WIDTH		8
 
	/************** Operation Code in instructions ****************/
	`define OP_NOP			4'b0000
	`define OP_ADD			4'b0001
	`define OP_SUB			4'b0010
	`define OP_AND			4'b0011
	`define OP_OR			4'b0100
	`define OP_XOR			4'b0101
	`define OP_SL			4'b0110
	`define OP_SR			4'b0111
	`define OP_SRU			4'b1000
	`define OP_ADDI			4'b1001
	`define OP_LD			4'b1010
	`define OP_ST			4'b1011
	`define OP_BZ			4'b1100
	
	/************** ALU operation command ****************/
	`define ALU_NC			3'bxxx		// not care
	`define ALU_ADD			3'b000
	`define ALU_SUB			3'b001
	`define ALU_AND			3'b010
	`define ALU_OR			3'b011
	`define ALU_XOR			3'b100
	`define ALU_SL			3'b101
	`define ALU_SR			3'b110
	`define ALU_SRU			3'b111
	
	/************** Branch condition code ****************/
	`define BRANCH_Z		3'b000
	//`define BRANCH_GT		3'b001
	//`define BRANCH_LE		3'b010
module mips_16_core_top
    (
        input						clk,
        input						rst,

        output	[`PC_WIDTH-1:0]		pc
    );
    wire 						pipeline_stall_n ;
    wire	[5:0]				branch_offset_imm;
    wire						branch_taken;
    wire	[15:0]				instruction;
    wire	[56:0]				ID_pipeline_reg_out;
    wire	[37:0]				EX_pipeline_reg_out;
    wire	[36:0]				MEM_pipeline_reg_out;

    wire	[2:0]				reg_read_addr_1;	// register file read port 1 address
    wire	[2:0]				reg_read_addr_2;	// register file read port 2 address
    wire	[15:0]				reg_read_data_1;	// register file read port 1 data
    wire	[15:0]				reg_read_data_2;	// register file read port 2 data
    wire	[2:0]				decoding_op_src1;		//source_1 register number
    wire	[2:0]				decoding_op_src2;		//source_2 register number
    wire	[2:0]				ex_op_dest;				//EX stage destinaton register number
    wire	[2:0]				mem_op_dest;			//MEM stage destinaton register number
    wire	[2:0]				wb_op_dest;				//WB stage destinaton register number
    wire						reg_write_en;
    wire	[2:0]				reg_write_dest;
    wire	[15:0]				reg_write_data;


    wire  IF_stage_inst_clk;
    wire  IF_stage_inst_rst;
    wire  IF_stage_inst_instruction_fetch_en;
    wire [5:0] IF_stage_inst_branch_offset_imm;
    wire  IF_stage_inst_branch_taken;
    reg [-1:0] IF_stage_inst_pc;
    wire [15:0] IF_stage_inst_instruction;
    assign IF_stage_inst_clk = clk;
    assign IF_stage_inst_rst = rst;
    assign IF_stage_inst_instruction_fetch_en = pipeline_stall_n;
    assign IF_stage_inst_branch_offset_imm = branch_offset_imm;
    assign IF_stage_inst_branch_taken = branch_taken;
    assign pc = IF_stage_inst_pc;
    assign instruction = IF_stage_inst_instruction;

    always @(  posedge   IF_stage_inst_clk or posedge  IF_stage_inst_rst )
    begin
        if ( IF_stage_inst_rst )
        begin
            IF_stage_inst_pc  <='b0;
        end
        else
        begin
            if ( IF_stage_inst_instruction_fetch_en )
            begin
                if ( IF_stage_inst_branch_taken )
                    IF_stage_inst_pc  <= IF_stage_inst_pc +{{(-6){ IF_stage_inst_branch_offset_imm [5]}}, IF_stage_inst_branch_offset_imm [5:0]};
                else
                    IF_stage_inst_pc  <= IF_stage_inst_pc +'d1;
            end
        end
    end


    wire  IF_stage_inst_imem_clk;
    wire [-1:0] IF_stage_inst_imem_pc;
    wire [15:0] IF_stage_inst_imem_instruction;
    assign IF_stage_inst_imem_clk = IF_stage_inst_clk;
    assign IF_stage_inst_imem_pc = IF_stage_inst_pc;
    assign IF_stage_inst_instruction = IF_stage_inst_imem_instruction;

    wire[-1:0] IF_stage_inst_imem_rom_addr = IF_stage_inst_imem_pc [-1:0];
    always @(*)
    case ( IF_stage_inst_imem_rom_addr )
        4 'b0000:
            IF_stage_inst_imem_instruction  =16'b1001001000001000;
        4 'b0001:
            IF_stage_inst_imem_instruction  =16'b1001010001001000;
        4 'b0010:
            IF_stage_inst_imem_instruction  =16'b1001011010001000;
        4 'b0011:
            IF_stage_inst_imem_instruction  =16'b0001100010011000;
        4 'b0100:
            IF_stage_inst_imem_instruction  =16'b1011100001000010;
        4 'b0101:
            IF_stage_inst_imem_instruction  =16'b1010101001000010;
        4 'b0110:
            IF_stage_inst_imem_instruction  =16'b0010110100101000;
        4 'b0111:
            IF_stage_inst_imem_instruction  =16'b1100000110111000;
        4 'b1000:
            IF_stage_inst_imem_instruction  =16'b1001111111000001;
        4 'b1001:
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
        4 'b1010:
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
        4 'b1011:
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
        4 'b1100:
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
        4 'b1101:
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
        4 'b1110:
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
        4 'b1111:
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
        default :
            IF_stage_inst_imem_instruction  =16'b0000000000000000;
    endcase





    wire  ID_stage_inst_clk;
    wire  ID_stage_inst_rst;
    wire  ID_stage_inst_instruction_decode_en;
    reg [56:
         0] ID_stage_inst_pipeline_reg_out;
    wire [15:
          0] ID_stage_inst_instruction;
    wire [5:
          0] ID_stage_inst_branch_offset_imm;
    reg  ID_stage_inst_branch_taken;
    wire [2:
          0] ID_stage_inst_reg_read_addr_1;
    wire [2:
          0] ID_stage_inst_reg_read_addr_2;
    wire [15:
          0] ID_stage_inst_reg_read_data_1;
    wire [15:
          0] ID_stage_inst_reg_read_data_2;
    wire [2:
          0] ID_stage_inst_decoding_op_src1;
    wire [2:
          0] ID_stage_inst_decoding_op_src2;
    assign ID_stage_inst_clk = clk;
    assign ID_stage_inst_rst = rst;
    assign ID_stage_inst_instruction_decode_en = pipeline_stall_n;
    assign ID_pipeline_reg_out = ID_stage_inst_pipeline_reg_out;
    assign ID_stage_inst_instruction = instruction;
    assign branch_offset_imm = ID_stage_inst_branch_offset_imm;
    assign branch_taken = ID_stage_inst_branch_taken;
    assign reg_read_addr_1 = ID_stage_inst_reg_read_addr_1;
    assign reg_read_addr_2 = ID_stage_inst_reg_read_addr_2;
    assign ID_stage_inst_reg_read_data_1 = reg_read_data_1;
    assign ID_stage_inst_reg_read_data_2 = reg_read_data_2;
    assign decoding_op_src1 = ID_stage_inst_decoding_op_src1;
    assign decoding_op_src2 = ID_stage_inst_decoding_op_src2;

    reg[15:
        0] ID_stage_inst_instruction_reg ;
    wire[3:
         0] ID_stage_inst_ir_op_code ;
    wire[2:
         0] ID_stage_inst_ir_dest ;
    wire[2:
         0] ID_stage_inst_ir_src1 ;
    wire[2:
         0] ID_stage_inst_ir_src2 ;
    wire[5:
         0] ID_stage_inst_ir_imm ;
    reg ID_stage_inst_write_back_en ;
    wire[2:
         0] ID_stage_inst_write_back_dest ;
    reg ID_stage_inst_write_back_result_mux ;
    wire ID_stage_inst_mem_write_en ;
    wire[15:
         0] ID_stage_inst_mem_write_data ;
    reg[2:
        0] ID_stage_inst_ex_alu_cmd ;
    wire[15:
         0] ID_stage_inst_ex_alu_src1 ;
    wire[15:
         0] ID_stage_inst_ex_alu_src2 ;
    reg ID_stage_inst_alu_src2_mux ;
    wire ID_stage_inst_decoding_op_is_branch ;
    wire ID_stage_inst_decoding_op_is_store ;
    wire[3:
         0] ID_stage_inst_ir_op_code_with_bubble ;
    wire[2:
         0] ID_stage_inst_ir_dest_with_bubble ;
    always @(  posedge   ID_stage_inst_clk or posedge  ID_stage_inst_rst )
    begin
        if ( ID_stage_inst_rst )
        begin
            ID_stage_inst_instruction_reg  <=0;
        end
        else
        begin
            if ( ID_stage_inst_instruction_decode_en )
            begin
                ID_stage_inst_instruction_reg  <= ID_stage_inst_instruction ;
            end
        end
    end

    assign  ID_stage_inst_ir_op_code = ID_stage_inst_instruction_reg [15:
            12];
    assign  ID_stage_inst_ir_dest = ID_stage_inst_instruction_reg [11:
            9];
    assign  ID_stage_inst_ir_src1 = ID_stage_inst_instruction_reg [8:
            6];
    assign  ID_stage_inst_ir_src2 =( ID_stage_inst_decoding_op_is_store )? ID_stage_inst_instruction_reg [11:9]: ID_stage_inst_instruction_reg [5:3];
    assign  ID_stage_inst_ir_imm = ID_stage_inst_instruction_reg [5:
            0];
    assign  ID_stage_inst_ir_op_code_with_bubble =( ID_stage_inst_instruction_decode_en )? ID_stage_inst_ir_op_code :0;
    assign  ID_stage_inst_ir_dest_with_bubble =( ID_stage_inst_instruction_decode_en )? ID_stage_inst_ir_dest :0;
    always @(*)
    begin
        if ( ID_stage_inst_rst )
        begin
            ID_stage_inst_write_back_en  =0;
            ID_stage_inst_write_back_result_mux  =0;
            ID_stage_inst_ex_alu_cmd  =0;
            ID_stage_inst_alu_src2_mux  =0;
        end
        else
        begin
            case( ID_stage_inst_ir_op_code_with_bubble )
                :
                begin
                    write_back_en=0;
                    write_back_result_mux=1'bx;
                    ex_alu_cmd=;
                    alu_src2_mux=1'bx;
                end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=0;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=0;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=0;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=0;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=1'bx;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=0;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=0;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=0;end:begin  write_back_en=1;  write_back_result_mux=0;  ex_alu_cmd=;  alu_src2_mux=1;end:begin  write_back_en=1;  write_back_result_mux=1;  ex_alu_cmd=;  alu_src2_mux=1;end:begin  write_back_en=0;  write_back_result_mux=1'bx;  ex_alu_cmd=;  alu_src2_mux=1;end:begin  write_back_en=0;  write_back_result_mux=1'bx;  ex_alu_cmd=;  alu_src2_mux=1;enddefault:begin  write_back_en=0;  write_back_result_mux=1'bx;  ex_alu_cmd=;  alu_src2_mux=1'bx;endendcaseendend
                        assign  ID_stage_inst_decoding_op_is_branch =( ID_stage_inst_ir_op_code ==)?1:0;
                        assign  ID_stage_inst_decoding_op_is_store =( ID_stage_inst_ir_op_code ==)?1:0;
                        assign  ID_stage_inst_mem_write_data = ID_stage_inst_reg_read_data_2 ;
                        assign  ID_stage_inst_mem_write_en = ID_stage_inst_decoding_op_is_store ;
                        assign  ID_stage_inst_write_back_dest = ID_stage_inst_ir_dest_with_bubble ;
                        assign  ID_stage_inst_ex_alu_src1 = ID_stage_inst_reg_read_data_1 ;
                        assign  ID_stage_inst_ex_alu_src2 =( ID_stage_inst_alu_src2_mux )?{{10{ ID_stage_inst_ir_imm [5]}}, ID_stage_inst_ir_imm }: ID_stage_inst_reg_read_data_2 ;
                        always @(  posedge   ID_stage_inst_clk or posedge  ID_stage_inst_rst )
                        begin
                            if ( ID_stage_inst_rst )
                            begin
                                ID_stage_inst_pipeline_reg_out  [56:0]<=0;
                            end
                            else
                            begin
                                ID_stage_inst_pipeline_reg_out  [56:0]<={ ID_stage_inst_ex_alu_cmd [2:0], ID_stage_inst_ex_alu_src1 [15:0], ID_stage_inst_ex_alu_src2 [15:0], ID_stage_inst_mem_write_en , ID_stage_inst_mem_write_data [15:0], ID_stage_inst_write_back_en , ID_stage_inst_write_back_dest [2:0], ID_stage_inst_write_back_result_mux };
                            end
                        end

                        assign  ID_stage_inst_reg_read_addr_1 = ID_stage_inst_ir_src1 ;
                        assign  ID_stage_inst_reg_read_addr_2 = ID_stage_inst_ir_src2 ;
                        always @(*)
                        begin
                            if ( ID_stage_inst_decoding_op_is_branch )
                            begin
                                case ( ID_stage_inst_ir_dest_with_bubble )
                                    :
                                    begin
                                        if ( ID_stage_inst_reg_read_data_1 ==0)
                                            ID_stage_inst_branch_taken  =1;
                                        else
                                            ID_stage_inst_branch_taken  =0;
                                    end
                                    default:
                                    begin
                                        ID_stage_inst_branch_taken  =0;
                                    end
                                endcase
                            end
                            else
                            begin
                                ID_stage_inst_branch_taken  =0;
                            end
                        end

                        assign  ID_stage_inst_branch_offset_imm = ID_stage_inst_ir_imm ;
                        assign  ID_stage_inst_decoding_op_src1 = ID_stage_inst_ir_src1 ;
                        assign  ID_stage_inst_decoding_op_src2 =( ID_stage_inst_ir_op_code <missing ')'>==||  ir_op_code==||  ir_op_code==||  ir_op_code==)?3'b000:  ir_src2;



                        wire  EX_stage_inst_clk;
                        wire  EX_stage_inst_rst;
                        wire [56:0] EX_stage_inst_pipeline_reg_in;
                            reg [37:0] EX_stage_inst_pipeline_reg_out;
                                wire [2:0] EX_stage_inst_ex_op_dest;
                                    assign EX_stage_inst_clk = clk;
                                    assign EX_stage_inst_rst = rst;
                                    assign EX_stage_inst_pipeline_reg_in = ID_pipeline_reg_out;
                                    assign EX_pipeline_reg_out = EX_stage_inst_pipeline_reg_out;
                                    assign ex_op_dest = EX_stage_inst_ex_op_dest;

                                    wire[2:0] EX_stage_inst_alu_cmd = EX_stage_inst_pipeline_reg_in [56:54];
                                            wire[15:0] EX_stage_inst_alu_src1 = EX_stage_inst_pipeline_reg_in [53:38];
                                                    wire[15:0] EX_stage_inst_alu_src2 = EX_stage_inst_pipeline_reg_in [37:22];
                                                            wire[15:0] EX_stage_inst_ex_alu_result ;

                                                                wire [15:0] EX_stage_inst_alu_inst_a;
                                                                    wire [15:0] EX_stage_inst_alu_inst_b;
                                                                        wire [2:0] EX_stage_inst_alu_inst_cmd;
                                                                            reg [15:0] EX_stage_inst_alu_inst_r;
                                                                                assign EX_stage_inst_alu_inst_a = EX_stage_inst_alu_src1;
                                                                                assign EX_stage_inst_alu_inst_b = EX_stage_inst_alu_src2;
                                                                                assign EX_stage_inst_alu_inst_cmd = EX_stage_inst_alu_cmd;
                                                                                assign EX_stage_inst_ex_alu_result = EX_stage_inst_alu_inst_r;

                                                                                always @(*)
                                                                                begin
                                                                                    case ( EX_stage_inst_alu_inst_cmd )
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  =
                                                                                            16 'bx;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  = EX_stage_inst_alu_inst_a + EX_stage_inst_alu_inst_b ;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  =
                                                                                            EX_stage_inst_alu_inst_a  - EX_stage_inst_alu_inst_b ;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  = EX_stage_inst_alu_inst_a & EX_stage_inst_alu_inst_b ;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  =
                                                                                            EX_stage_inst_alu_inst_a  | EX_stage_inst_alu_inst_b ;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  = EX_stage_inst_alu_inst_a ^ EX_stage_inst_alu_inst_b ;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  =
                                                                                            EX_stage_inst_alu_inst_a  << EX_stage_inst_alu_inst_b ;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  ={{16{ EX_stage_inst_alu_inst_a [15]}}, EX_stage_inst_alu_inst_a }>> EX_stage_inst_alu_inst_b ;
                                                                                        :
                                                                                            EX_stage_inst_alu_inst_r  =
                                                                                            { 16'b0, EX_stage_inst_alu_inst_a }>> EX_stage_inst_alu_inst_b ;
                                                                                        default :
                                                                                        begin
                                                                                            EX_stage_inst_alu_inst_r  =0;
                                                                                        end
                                                                                    endcase
                                                                                end


                        always @( posedge  EX_stage_inst_clk )
                        begin
                            if ( EX_stage_inst_rst )
                            begin
                                EX_stage_inst_pipeline_reg_out  [37:0]<=0;
                            end
                            else
                            begin
                                EX_stage_inst_pipeline_reg_out  [37:22]<= EX_stage_inst_ex_alu_result ;
                                EX_stage_inst_pipeline_reg_out  [21:0]<= EX_stage_inst_pipeline_reg_in [21:0];
                            end
                        end

                        assign  EX_stage_inst_ex_op_dest = EX_stage_inst_pipeline_reg_in [3:1];



                            wire  MEM_stage_inst_clk;
                            wire  MEM_stage_inst_rst;
                            wire [37:0] MEM_stage_inst_pipeline_reg_in;
                                reg [36:0] MEM_stage_inst_pipeline_reg_out;
                                    wire [2:0] MEM_stage_inst_mem_op_dest;
                                        assign MEM_stage_inst_clk = clk;
                                        assign MEM_stage_inst_rst = rst;
                                        assign MEM_stage_inst_pipeline_reg_in = EX_pipeline_reg_out;
                                        assign MEM_pipeline_reg_out = MEM_stage_inst_pipeline_reg_out;
                                        assign mem_op_dest = MEM_stage_inst_mem_op_dest;

                                        wire[15:0] MEM_stage_inst_ex_alu_result = MEM_stage_inst_pipeline_reg_in [37:22];
                                                wire MEM_stage_inst_mem_write_en = MEM_stage_inst_pipeline_reg_in [21];
                                                wire[15:0] MEM_stage_inst_mem_write_data = MEM_stage_inst_pipeline_reg_in [20:5];
                                                        wire[15:0] MEM_stage_inst_mem_read_data ;

                                                            wire  MEM_stage_inst_dmem_clk;
                                                            wire [15:0] MEM_stage_inst_dmem_mem_access_addr;
                                                                wire [15:0] MEM_stage_inst_dmem_mem_write_data;
                                                                    wire  MEM_stage_inst_dmem_mem_write_en;
                                                                    wire [15:0] MEM_stage_inst_dmem_mem_read_data;
                                                                        assign MEM_stage_inst_dmem_clk = MEM_stage_inst_clk;
                                                                        assign MEM_stage_inst_dmem_mem_access_addr = MEM_stage_inst_ex_alu_result;
                                                                        assign MEM_stage_inst_dmem_mem_write_data = MEM_stage_inst_mem_write_data;
                                                                        assign MEM_stage_inst_dmem_mem_write_en = MEM_stage_inst_mem_write_en;
                                                                        assign MEM_stage_inst_mem_read_data = MEM_stage_inst_dmem_mem_read_data;

                                                                        reg[15:0] MEM_stage_inst_dmem_ram [(2**) -1:0];
                                                                                wire[-1:0] MEM_stage_inst_dmem_ram_addr = MEM_stage_inst_dmem_mem_access_addr [-1:0];
                                                                                        always @( posedge  MEM_stage_inst_dmem_clk )
                                                                                            if ( MEM_stage_inst_dmem_mem_write_en )
                                                                                            MEM_stage_inst_dmem_ram  [ MEM_stage_inst_dmem_ram_addr ]<= MEM_stage_inst_dmem_mem_write_data ;

                                                                                            assign  MEM_stage_inst_dmem_mem_read_data = MEM_stage_inst_dmem_ram [ MEM_stage_inst_dmem_ram_addr ];

                                                                                            always @( posedge  MEM_stage_inst_clk )
                                                                                            begin
                                                                                                if ( MEM_stage_inst_rst )
                                                                                                    begin
                                                                                                        MEM_stage_inst_pipeline_reg_out  [36:0]<=0;
                                                                                                    end
                                                                                                    else
                                                                                                    begin
                                                                                                        MEM_stage_inst_pipeline_reg_out  [36:21]<= MEM_stage_inst_ex_alu_result ;
                                                                                                        MEM_stage_inst_pipeline_reg_out  [20:5]<= MEM_stage_inst_mem_read_data ;
                                                                                                        MEM_stage_inst_pipeline_reg_out  [4:0]<= MEM_stage_inst_pipeline_reg_in [4:0];
                                                                                                    end
                                                                                                end

                        assign  MEM_stage_inst_mem_op_dest = MEM_stage_inst_pipeline_reg_in [3:1];



                            wire [36:0] WB_stage_inst_pipeline_reg_in;
                                wire  WB_stage_inst_reg_write_en;
                                wire [2:0] WB_stage_inst_reg_write_dest;
                                    wire [15:0] WB_stage_inst_reg_write_data;
                                        wire [2:0] WB_stage_inst_wb_op_dest;
                                            assign WB_stage_inst_pipeline_reg_in = MEM_pipeline_reg_out;
                                            assign reg_write_en = WB_stage_inst_reg_write_en;
                                            assign reg_write_dest = WB_stage_inst_reg_write_dest;
                                            assign reg_write_data = WB_stage_inst_reg_write_data;
                                            assign wb_op_dest = WB_stage_inst_wb_op_dest;

                                            wire[15:0] WB_stage_inst_ex_alu_result = WB_stage_inst_pipeline_reg_in [36:21];
                                                    wire[15:0] WB_stage_inst_mem_read_data = WB_stage_inst_pipeline_reg_in [20:5];
                                                            wire WB_stage_inst_write_back_en = WB_stage_inst_pipeline_reg_in [4];
                                                            wire[2:0] WB_stage_inst_write_back_dest = WB_stage_inst_pipeline_reg_in [3:1];
                                                                    wire WB_stage_inst_write_back_result_mux = WB_stage_inst_pipeline_reg_in [0];
                                                                    assign  WB_stage_inst_reg_write_en = WB_stage_inst_write_back_en ;
                                                                    assign  WB_stage_inst_reg_write_dest = WB_stage_inst_write_back_dest ;
                                                                    assign  WB_stage_inst_reg_write_data =( WB_stage_inst_write_back_result_mux )? WB_stage_inst_mem_read_data : WB_stage_inst_ex_alu_result ;
                                                                    assign  WB_stage_inst_wb_op_dest = WB_stage_inst_pipeline_reg_in [3:1];



                                                                        wire  register_file_inst_clk;
                                                                        wire  register_file_inst_rst;
                                                                        wire  register_file_inst_reg_write_en;
                                                                        wire [2:0] register_file_inst_reg_write_dest;
                                                                            wire [15:0] register_file_inst_reg_write_data;
                                                                                wire [2:0] register_file_inst_reg_read_addr_1;
                                                                                    wire [15:0] register_file_inst_reg_read_data_1;
                                                                                        wire [2:0] register_file_inst_reg_read_addr_2;
                                                                                            wire [15:0] register_file_inst_reg_read_data_2;
                                                                                                assign register_file_inst_clk = clk;
                                                                                                assign register_file_inst_rst = rst;
                                                                                                assign register_file_inst_reg_write_en = reg_write_en;
                                                                                                assign register_file_inst_reg_write_dest = reg_write_dest;
                                                                                                assign register_file_inst_reg_write_data = reg_write_data;
                                                                                                assign register_file_inst_reg_read_addr_1 = reg_read_addr_1;
                                                                                                assign reg_read_data_1 = register_file_inst_reg_read_data_1;
                                                                                                assign register_file_inst_reg_read_addr_2 = reg_read_addr_2;
                                                                                                assign reg_read_data_2 = register_file_inst_reg_read_data_2;

                                                                                                reg[15:0] register_file_inst_reg_array [7:0];
                                                                                                        always @(  posedge   register_file_inst_clk or posedge  register_file_inst_rst )
                                                                                                        begin
                                                                                                            if ( register_file_inst_rst )
                                                                                                            begin
                                                                                                                register_file_inst_reg_array  [0]<=15'b0;
                                                                                                                register_file_inst_reg_array  [1]<=15'b0;
                                                                                                                register_file_inst_reg_array  [2]<=15'b0;
                                                                                                                register_file_inst_reg_array  [3]<=15'b0;
                                                                                                                register_file_inst_reg_array  [4]<=15'b0;
                                                                                                                register_file_inst_reg_array  [5]<=15'b0;
                                                                                                                register_file_inst_reg_array  [6]<=15'b0;
                                                                                                                register_file_inst_reg_array  [7]<=15'b0;
                                                                                                            end
                                                                                                            else
                                                                                                            begin
                                                                                                                if ( register_file_inst_reg_write_en )
                                                                                                                begin
                                                                                                                    register_file_inst_reg_array  [ register_file_inst_reg_write_dest ]<= register_file_inst_reg_write_data ;
                                                                                                                end
                                                                                                            end
                                                                                                        end

                        assign  register_file_inst_reg_read_data_1 =( register_file_inst_reg_read_addr_1 ==0)?15'b0: register_file_inst_reg_array [ register_file_inst_reg_read_addr_1 ];
                        assign  register_file_inst_reg_read_data_2 =( register_file_inst_reg_read_addr_2 ==0)?15'b0: register_file_inst_reg_array [ register_file_inst_reg_read_addr_2 ];



                        wire [2:0] hazard_detection_unit_inst_decoding_op_src1;
                            wire [2:0] hazard_detection_unit_inst_decoding_op_src2;
                                wire [2:0] hazard_detection_unit_inst_ex_op_dest;
                                    wire [2:0] hazard_detection_unit_inst_mem_op_dest;
                                        wire [2:0] hazard_detection_unit_inst_wb_op_dest;
                                            reg  hazard_detection_unit_inst_pipeline_stall_n;
                                            assign hazard_detection_unit_inst_decoding_op_src1 = decoding_op_src1;
                                            assign hazard_detection_unit_inst_decoding_op_src2 = decoding_op_src2;
                                            assign hazard_detection_unit_inst_ex_op_dest = ex_op_dest;
                                            assign hazard_detection_unit_inst_mem_op_dest = mem_op_dest;
                                            assign hazard_detection_unit_inst_wb_op_dest = wb_op_dest;
                                            assign pipeline_stall_n = hazard_detection_unit_inst_pipeline_stall_n;

                                            always @(*)
                                            begin
                                                hazard_detection_unit_inst_pipeline_stall_n  =1;
                                                if ( hazard_detection_unit_inst_decoding_op_src1 !=0&&( hazard_detection_unit_inst_decoding_op_src1 == hazard_detection_unit_inst_ex_op_dest || hazard_detection_unit_inst_decoding_op_src1 == hazard_detection_unit_inst_mem_op_dest || hazard_detection_unit_inst_decoding_op_src1 == hazard_detection_unit_inst_wb_op_dest ))
                                                    hazard_detection_unit_inst_pipeline_stall_n  =0;
                                                if ( hazard_detection_unit_inst_decoding_op_src2 !=0&&( hazard_detection_unit_inst_decoding_op_src2 == hazard_detection_unit_inst_ex_op_dest || hazard_detection_unit_inst_decoding_op_src2 == hazard_detection_unit_inst_mem_op_dest || hazard_detection_unit_inst_decoding_op_src2 == hazard_detection_unit_inst_wb_op_dest ))
                                                    hazard_detection_unit_inst_pipeline_stall_n  =0;
                                            end



                    endmodule
